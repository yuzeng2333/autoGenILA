module SDP_Y_CORE_Y_mul_core(nvdla_core_clk, nvdla_core_rstn, chn_mul_in_rsc_z, chn_mul_in_rsc_vz, chn_mul_in_rsc_lz, chn_mul_op_rsc_z, chn_mul_op_rsc_vz, chn_mul_op_rsc_lz, cfg_mul_bypass_rsc_triosy_lz, cfg_mul_prelu_rsc_triosy_lz, cfg_mul_src_rsc_triosy_lz, cfg_mul_op_rsc_triosy_lz, cfg_truncate_rsc_triosy_lz, cfg_precision, chn_mul_out_rsc_z, chn_mul_out_rsc_vz, chn_mul_out_rsc_lz, chn_mul_in_rsci_oswt, chn_mul_in_rsci_oswt_unreg, chn_mul_op_rsci_oswt, chn_mul_op_rsci_oswt_unreg, cfg_mul_bypass_rsci_d, cfg_mul_prelu_rsci_d, cfg_mul_src_rsci_d, cfg_mul_op_rsci_d, cfg_truncate_rsci_d, chn_mul_out_rsci_oswt, chn_mul_out_rsci_oswt_unreg, cfg_mul_bypass_rsc_triosy_obj_oswt, cfg_mul_prelu_rsc_triosy_obj_oswt, cfg_mul_src_rsc_triosy_obj_oswt, cfg_mul_op_rsc_triosy_obj_oswt, cfg_truncate_rsc_triosy_obj_oswt, cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_pff);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10010" *)
  wire _00000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10010" *)
  wire _00001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10010" *)
  wire _00002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10027" *)
  wire [21:0] _00003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10027" *)
  wire [21:0] _00004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10027" *)
  wire [21:0] _00005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10027" *)
  wire [21:0] _00006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10027" *)
  wire [21:0] _00007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10027" *)
  wire [21:0] _00008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10027" *)
  wire [21:0] _00009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10027" *)
  wire [21:0] _00010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10044" *)
  wire [22:0] _00022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10146" *)
  wire [7:0] _00023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10146" *)
  wire [7:0] _00024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10146" *)
  wire [7:0] _00025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10146" *)
  wire [7:0] _00026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10146" *)
  wire [7:0] _00027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10146" *)
  wire [7:0] _00028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10146" *)
  wire [7:0] _00029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10146" *)
  wire [7:0] _00030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8544" *)
  wire _00031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7931" *)
  wire _00032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8609" *)
  wire _00033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8068" *)
  wire _00034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8674" *)
  wire _00035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8205" *)
  wire _00036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8739" *)
  wire _00037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8342" *)
  wire _00038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8609" *)
  wire _00039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8018" *)
  wire _00040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8674" *)
  wire _00041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8155" *)
  wire _00042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8739" *)
  wire _00043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8292" *)
  wire _00044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8544" *)
  wire _00045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7881" *)
  wire _00046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8588" *)
  wire _00047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7978" *)
  wire _00048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8653" *)
  wire _00049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8115" *)
  wire _00050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8718" *)
  wire _00051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8252" *)
  wire _00052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8523" *)
  wire _00053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7841" *)
  wire _00054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8503" *)
  wire _00055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7828" *)
  wire _00056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8568" *)
  wire _00057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7965" *)
  wire _00058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8633" *)
  wire _00059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8102" *)
  wire _00060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8698" *)
  wire _00061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8239" *)
  wire _00062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8847" *)
  wire _00063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8325" *)
  wire _00064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9027" *)
  wire _00065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7715" *)
  wire _00066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8315" *)
  wire _00067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8763" *)
  wire _00068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7914" *)
  wire _00069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8979" *)
  wire _00070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7559" *)
  wire _00071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7904" *)
  wire _00072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8791" *)
  wire _00073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8051" *)
  wire _00074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8995" *)
  wire _00075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7611" *)
  wire _00076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8041" *)
  wire _00077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8819" *)
  wire _00078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8188" *)
  wire _00079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9011" *)
  wire _00080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7663" *)
  wire _00081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8178" *)
  wire _00082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8780" *)
  wire _00083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7776" *)
  wire _00084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8808" *)
  wire _00085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7786" *)
  wire _00086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8836" *)
  wire _00087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7796" *)
  wire _00088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8864" *)
  wire _00089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7806" *)
  wire _00090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8523" *)
  wire [7:0] _00091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7816" *)
  wire [7:0] _00092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8588" *)
  wire [7:0] _00093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7953" *)
  wire [7:0] _00094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8653" *)
  wire [7:0] _00095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8090" *)
  wire [7:0] _00096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8718" *)
  wire [7:0] _00097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8227" *)
  wire [7:0] _00098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8875" *)
  wire [47:0] _00099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8907" *)
  wire [47:0] _00100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8928" *)
  wire [47:0] _00101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8949" *)
  wire [47:0] _00102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7776" *)
  wire [31:0] _00103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7871" *)
  wire _00104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7786" *)
  wire [31:0] _00105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8008" *)
  wire _00106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7796" *)
  wire [31:0] _00107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8145" *)
  wire _00108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7806" *)
  wire [31:0] _00109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8282" *)
  wire _00110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8771" *)
  wire _00111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7871" *)
  wire _00112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8799" *)
  wire _00113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8008" *)
  wire _00114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8827" *)
  wire _00115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8145" *)
  wire _00116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8855" *)
  wire _00117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8282" *)
  wire _00118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8386" *)
  wire _00119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7501" *)
  wire _00120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7750" *)
  wire _00121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9035" *)
  wire _00122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8414" *)
  wire _00123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7537" *)
  wire _00124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7904" *)
  wire _00125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8386" *)
  wire _00126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7501" *)
  wire _00127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7750" *)
  wire _00128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9045" *)
  wire _00129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8443" *)
  wire _00130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7589" *)
  wire _00131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8041" *)
  wire _00132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8386" *)
  wire _00133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7501" *)
  wire _00134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7750" *)
  wire _00135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9055" *)
  wire _00136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8455" *)
  wire _00137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7641" *)
  wire _00138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8178" *)
  wire _00139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8386" *)
  wire _00140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7501" *)
  wire _00141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7750" *)
  wire _00142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9065" *)
  wire _00143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8467" *)
  wire _00144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7693" *)
  wire _00145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8315" *)
  wire _00146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8971" *)
  wire _00147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7527" *)
  wire _00148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8987" *)
  wire _00149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7579" *)
  wire _00150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9003" *)
  wire _00151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7631" *)
  wire _00152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9019" *)
  wire _00153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7683" *)
  wire _00154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9035" *)
  wire _00155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8414" *)
  wire _00156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7493" *)
  wire _00157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9045" *)
  wire _00158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8443" *)
  wire _00159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7571" *)
  wire _00160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9055" *)
  wire _00161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8455" *)
  wire _00162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7623" *)
  wire _00163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9065" *)
  wire _00164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8467" *)
  wire _00165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7675" *)
  wire _00166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7501" *)
  wire [127:0] _00167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7750" *)
  wire [127:0] _00168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8386" *)
  wire [127:0] _00169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8426" *)
  wire [31:0] _00170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8435" *)
  wire _00171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9075" *)
  wire _00172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8493" *)
  wire _00173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8386" *)
  wire [9:0] _00174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8897" *)
  wire [9:0] _00175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7379" *)
  wire _00176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7393" *)
  wire _00177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7379" *)
  wire _00178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7477" *)
  wire _00179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7431" *)
  wire [21:0] _00181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7431" *)
  wire [7:0] _00182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7431" *)
  wire [21:0] _00184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7431" *)
  wire [7:0] _00185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7431" *)
  wire [21:0] _00188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7431" *)
  wire [7:0] _00189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7431" *)
  wire [21:0] _00192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7431" *)
  wire [7:0] _00193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7379" *)
  wire _00196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7537" *)
  wire [30:0] _00197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7589" *)
  wire [30:0] _00198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7641" *)
  wire [30:0] _00199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7693" *)
  wire [30:0] _00200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8544" *)
  wire [22:0] _00201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7892" *)
  wire [22:0] _00202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8535" *)
  wire [7:0] _00203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8609" *)
  wire [22:0] _00204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8029" *)
  wire [22:0] _00205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8600" *)
  wire [7:0] _00206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8674" *)
  wire [22:0] _00207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8166" *)
  wire [22:0] _00208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8665" *)
  wire [7:0] _00209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8739" *)
  wire [22:0] _00210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8303" *)
  wire [22:0] _00211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8730" *)
  wire [7:0] _00212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7750" *)
  wire _00213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8386" *)
  wire _00214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7501" *)
  wire _00215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8378" *)
  wire _00216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7485" *)
  wire _00217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7741" *)
  wire _00218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7881" *)
  wire _00219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8544" *)
  wire _00220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7922" *)
  wire _00221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8513" *)
  wire [22:0] _00222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8523" *)
  wire _00223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7851" *)
  wire _00224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9083" *)
  wire _00225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8885" *)
  wire _00226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7547" *)
  wire _00227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7861" *)
  wire _00228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9093" *)
  wire [63:0] _00229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7559" *)
  wire [63:0] _00230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8558" *)
  wire _00231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7941" *)
  wire _00232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8558" *)
  wire _00233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7941" *)
  wire _00234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8018" *)
  wire _00235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8609" *)
  wire _00236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8059" *)
  wire _00237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8578" *)
  wire [22:0] _00238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8588" *)
  wire _00239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7988" *)
  wire _00240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9102" *)
  wire _00241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8916" *)
  wire _00242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7599" *)
  wire _00243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7998" *)
  wire _00244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9112" *)
  wire [63:0] _00245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7611" *)
  wire [63:0] _00246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8623" *)
  wire _00247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8078" *)
  wire _00248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8623" *)
  wire _00249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8078" *)
  wire _00250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8155" *)
  wire _00251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8674" *)
  wire _00252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8196" *)
  wire _00253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8643" *)
  wire [22:0] _00254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8653" *)
  wire _00255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8125" *)
  wire _00256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9121" *)
  wire _00257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8937" *)
  wire _00258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7651" *)
  wire _00259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8135" *)
  wire _00260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9131" *)
  wire [63:0] _00261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7663" *)
  wire [63:0] _00262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8688" *)
  wire _00263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8215" *)
  wire _00264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8688" *)
  wire _00265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8215" *)
  wire _00266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8292" *)
  wire _00267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8739" *)
  wire _00268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8333" *)
  wire _00269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8708" *)
  wire [22:0] _00270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8718" *)
  wire _00271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8262" *)
  wire _00272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9140" *)
  wire _00273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8959" *)
  wire _00274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7703" *)
  wire _00275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8272" *)
  wire _00276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9150" *)
  wire [63:0] _00277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7715" *)
  wire [63:0] _00278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8753" *)
  wire _00279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8352" *)
  wire _00280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8753" *)
  wire _00281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8352" *)
  wire _00282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8386" *)
  wire _00283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7501" *)
  wire _00284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7750" *)
  wire _00285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8479" *)
  wire _00286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7727" *)
  wire _00287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8364" *)
  wire _00288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8386" *)
  wire _00289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7501" *)
  wire _00290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7750" *)
  wire _00291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8479" *)
  wire _00292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7727" *)
  wire _00293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8364" *)
  wire _00294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8386" *)
  wire _00295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7501" *)
  wire _00296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7750" *)
  wire _00297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8479" *)
  wire _00298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7727" *)
  wire _00299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8364" *)
  wire _00300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8386" *)
  wire _00301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7501" *)
  wire _00302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7750" *)
  wire _00303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8479" *)
  wire _00304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7727" *)
  wire _00305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8364" *)
  wire _00306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7379" *)
  wire _00307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7469" *)
  wire _00308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7401" *)
  wire _00316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7527" *)
  wire _00317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7547" *)
  wire _00318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7559" *)
  wire _00319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7579" *)
  wire _00320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7599" *)
  wire _00321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7611" *)
  wire _00322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7631" *)
  wire _00323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7651" *)
  wire _00324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7663" *)
  wire _00325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7683" *)
  wire _00326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7703" *)
  wire _00327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7715" *)
  wire _00328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7828" *)
  wire _00329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7841" *)
  wire _00330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7851" *)
  wire _00331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7881" *)
  wire _00332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7931" *)
  wire _00333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7941" *)
  wire _00334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7941" *)
  wire _00335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7965" *)
  wire _00336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7978" *)
  wire _00337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7988" *)
  wire _00338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8018" *)
  wire _00339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8068" *)
  wire _00340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8078" *)
  wire _00341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8078" *)
  wire _00342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8102" *)
  wire _00343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8115" *)
  wire _00344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8125" *)
  wire _00345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8155" *)
  wire _00346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8205" *)
  wire _00347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8215" *)
  wire _00348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8215" *)
  wire _00349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8239" *)
  wire _00350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8252" *)
  wire _00351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8262" *)
  wire _00352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8292" *)
  wire _00353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8342" *)
  wire _00354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8352" *)
  wire _00355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8352" *)
  wire _00356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8414" *)
  wire _00357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8414" *)
  wire _00358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8443" *)
  wire _00359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8443" *)
  wire _00360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8455" *)
  wire _00361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8455" *)
  wire _00362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8467" *)
  wire _00363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8467" *)
  wire _00364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8493" *)
  wire _00365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8885" *)
  wire _00366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8916" *)
  wire _00367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8937" *)
  wire _00368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8959" *)
  wire _00369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7559" *)
  wire [63:0] _00370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7611" *)
  wire [63:0] _00371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7663" *)
  wire [63:0] _00372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7715" *)
  wire [63:0] _00373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *)
  wire [7:0] _00374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *)
  wire [7:0] _00375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *)
  wire [7:0] _00376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *)
  wire [7:0] _00377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *)
  wire [7:0] _00378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *)
  wire [7:0] _00379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *)
  wire [7:0] _00380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *)
  wire [7:0] _00381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _00382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _00383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _00384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _00385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _00386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _00387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _00388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _00389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _00390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _00391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _00392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _00393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _00394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _00395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _00396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _00397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _00398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _00399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _00400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _00401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _00402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _00403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _00404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _00405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4344" *)
  wire _00406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4344" *)
  wire _00407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4347" *)
  wire _00408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4349" *)
  wire _00409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4351" *)
  wire _00410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4353" *)
  wire _00411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4359" *)
  wire _00412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4371" *)
  wire _00413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4405" *)
  wire _00414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4410" *)
  wire _00415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4424" *)
  wire _00416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4443" *)
  wire _00417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4481" *)
  wire _00418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4494" *)
  wire _00419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *)
  wire _00420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *)
  wire _00421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *)
  wire _00422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *)
  wire _00423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4571" *)
  wire _00424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4575" *)
  wire _00425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4599" *)
  wire _00426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4603" *)
  wire _00427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4627" *)
  wire _00428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4631" *)
  wire _00429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4655" *)
  wire _00430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4659" *)
  wire _00431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4869" *)
  wire _00432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4871" *)
  wire _00433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4889" *)
  wire _00434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4891" *)
  wire _00435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4907" *)
  wire _00436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4909" *)
  wire _00437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4925" *)
  wire _00438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4927" *)
  wire _00439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4977" *)
  wire _00440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4977" *)
  wire _00441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4977" *)
  wire _00442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4978" *)
  wire _00443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4978" *)
  wire _00444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4978" *)
  wire _00445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4980" *)
  wire _00446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4980" *)
  wire _00447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7088" *)
  wire _00448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7091" *)
  wire _00449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7094" *)
  wire _00450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7097" *)
  wire _00451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7100" *)
  wire _00452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7100" *)
  wire _00453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7100" *)
  wire _00454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7101" *)
  wire _00455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7101" *)
  wire _00456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7101" *)
  wire _00457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7180" *)
  wire _00458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7271" *)
  wire _00459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7306" *)
  wire _00460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7309" *)
  wire _00461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7319" *)
  wire _00462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7359" *)
  wire _00463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7367" *)
  wire _00464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7371" *)
  wire _00465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7372" *)
  wire _00466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7373" *)
  wire _00467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7374" *)
  wire _00468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7387" *)
  wire _00469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7397" *)
  wire _00470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7473" *)
  wire _00471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7481" *)
  wire _00472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7489" *)
  wire _00473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7497" *)
  wire _00474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7532" *)
  wire _00475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7553" *)
  wire _00476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7575" *)
  wire _00477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7584" *)
  wire _00478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7605" *)
  wire _00479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7627" *)
  wire _00480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7636" *)
  wire _00481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7657" *)
  wire _00482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7679" *)
  wire _00483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7688" *)
  wire _00484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7709" *)
  wire _00485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7745" *)
  wire _00486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7820" *)
  wire _00487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7821" *)
  wire _00488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7834" *)
  wire _00489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7846" *)
  wire _00490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7856" *)
  wire _00491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7866" *)
  wire _00492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7897" *)
  wire _00493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7918" *)
  wire _00494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7927" *)
  wire _00495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7936" *)
  wire _00496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7957" *)
  wire _00497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7958" *)
  wire _00498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7971" *)
  wire _00499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7983" *)
  wire _00500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7993" *)
  wire _00501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8003" *)
  wire _00502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8034" *)
  wire _00503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8055" *)
  wire _00504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8064" *)
  wire _00505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8073" *)
  wire _00506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8094" *)
  wire _00507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8095" *)
  wire _00508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8108" *)
  wire _00509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8120" *)
  wire _00510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8130" *)
  wire _00511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8140" *)
  wire _00512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8171" *)
  wire _00513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8192" *)
  wire _00514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8201" *)
  wire _00515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8210" *)
  wire _00516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8231" *)
  wire _00517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8232" *)
  wire _00518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8245" *)
  wire _00519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8257" *)
  wire _00520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8267" *)
  wire _00521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8277" *)
  wire _00522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8308" *)
  wire _00523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8329" *)
  wire _00524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8338" *)
  wire _00525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8347" *)
  wire _00526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8382" *)
  wire _00527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8431" *)
  wire _00528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8439" *)
  wire _00529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8497" *)
  wire _00530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8498" *)
  wire _00531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8508" *)
  wire _00532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8518" *)
  wire _00533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8540" *)
  wire _00534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8573" *)
  wire _00535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8583" *)
  wire _00536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8605" *)
  wire _00537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8638" *)
  wire _00538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8648" *)
  wire _00539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8670" *)
  wire _00540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8703" *)
  wire _00541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8713" *)
  wire _00542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8735" *)
  wire _00543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8767" *)
  wire _00544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8768" *)
  wire _00545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8776" *)
  wire _00546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8785" *)
  wire _00547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8785" *)
  wire _00548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8795" *)
  wire _00549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8796" *)
  wire _00550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8804" *)
  wire _00551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8813" *)
  wire _00552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8813" *)
  wire _00553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8823" *)
  wire _00554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8824" *)
  wire _00555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8832" *)
  wire _00556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8841" *)
  wire _00557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8841" *)
  wire _00558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8851" *)
  wire _00559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8852" *)
  wire _00560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8860" *)
  wire _00561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8869" *)
  wire _00562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8869" *)
  wire _00563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8880" *)
  wire _00564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8881" *)
  wire _00565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8890" *)
  wire _00566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8890" *)
  wire _00567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8891" *)
  wire _00568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8902" *)
  wire _00569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8902" *)
  wire _00570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8902" *)
  wire _00571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8903" *)
  wire _00572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8911" *)
  wire _00573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8912" *)
  wire _00574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8921" *)
  wire _00575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8921" *)
  wire _00576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8922" *)
  wire _00577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8932" *)
  wire _00578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8933" *)
  wire _00579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8942" *)
  wire _00580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8942" *)
  wire _00581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8943" *)
  wire _00582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8954" *)
  wire _00583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8955" *)
  wire _00584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8964" *)
  wire _00585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8964" *)
  wire _00586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8965" *)
  wire _00587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8975" *)
  wire _00588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8975" *)
  wire _00589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8983" *)
  wire _00590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8991" *)
  wire _00591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8991" *)
  wire _00592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8999" *)
  wire _00593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9007" *)
  wire _00594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9007" *)
  wire _00595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9015" *)
  wire _00596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9023" *)
  wire _00597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9023" *)
  wire _00598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9031" *)
  wire _00599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9079" *)
  wire _00600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9089" *)
  wire _00601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9098" *)
  wire _00602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9108" *)
  wire _00603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9117" *)
  wire _00604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9127" *)
  wire _00605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9136" *)
  wire _00606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9146" *)
  wire _00607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9155" *)
  wire _00608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9235" *)
  wire _00609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9236" *)
  wire _00610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9254" *)
  wire _00611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9254" *)
  wire _00612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9272" *)
  wire _00613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9272" *)
  wire _00614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9289" *)
  wire _00615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9290" *)
  wire _00616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9331" *)
  wire _00617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9343" *)
  wire _00618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9357" *)
  wire _00619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9375" *)
  wire _00620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9393" *)
  wire _00621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9435" *)
  wire _00622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9444" *)
  wire _00623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9444" *)
  wire _00624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9447" *)
  wire _00625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9461" *)
  wire _00626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9497" *)
  wire _00627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9540" *)
  wire _00628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9549" *)
  wire _00629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9549" *)
  wire _00630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9552" *)
  wire _00631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9566" *)
  wire _00632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9602" *)
  wire _00633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9645" *)
  wire _00634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9654" *)
  wire _00635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9654" *)
  wire _00636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9657" *)
  wire _00637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9671" *)
  wire _00638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9708" *)
  wire _00639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9813" *)
  wire _00640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9831" *)
  wire _00641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9849" *)
  wire _00642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9867" *)
  wire _00643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9935" *)
  wire _00644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9935" *)
  wire _00645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9935" *)
  wire _00646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9935" *)
  wire _00647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *)
  wire _00648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *)
  wire _00649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *)
  wire _00650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *)
  wire _00651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *)
  wire _00652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *)
  wire _00653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *)
  wire _00654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *)
  wire _00655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9948" *)
  wire [21:0] _00656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9948" *)
  wire [21:0] _00657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9948" *)
  wire [21:0] _00658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9948" *)
  wire [21:0] _00659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *)
  wire [21:0] _00660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *)
  wire [21:0] _00661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *)
  wire [21:0] _00662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *)
  wire [21:0] _00663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *)
  wire [21:0] _00664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *)
  wire [21:0] _00665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *)
  wire [21:0] _00666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *)
  wire [21:0] _00667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9961" *)
  wire [22:0] _00668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9961" *)
  wire [22:0] _00669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9961" *)
  wire [22:0] _00670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9961" *)
  wire [22:0] _00671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *)
  wire [22:0] _00672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *)
  wire [22:0] _00673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *)
  wire [22:0] _00674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *)
  wire [22:0] _00675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *)
  wire [22:0] _00676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *)
  wire [22:0] _00677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *)
  wire [22:0] _00678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *)
  wire [22:0] _00679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9975" *)
  wire [22:0] _00680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9975" *)
  wire [22:0] _00681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9975" *)
  wire [22:0] _00682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9975" *)
  wire [22:0] _00683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *)
  wire [22:0] _00684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *)
  wire [22:0] _00685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *)
  wire [22:0] _00686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *)
  wire [22:0] _00687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *)
  wire [22:0] _00688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *)
  wire [22:0] _00689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *)
  wire [22:0] _00690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *)
  wire [22:0] _00691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *)
  wire [22:0] _00692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *)
  wire [22:0] _00693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *)
  wire [22:0] _00694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *)
  wire [22:0] _00695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9989" *)
  wire [7:0] _00696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9989" *)
  wire [7:0] _00697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9989" *)
  wire [7:0] _00698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9989" *)
  wire [7:0] _00699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *)
  wire [7:0] _00700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *)
  wire [7:0] _00701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *)
  wire [7:0] _00702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *)
  wire [7:0] _00703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *)
  wire [7:0] _00704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *)
  wire [7:0] _00705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *)
  wire [7:0] _00706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *)
  wire [7:0] _00707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4573" *)
  wire _00708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4590" *)
  wire _00709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4601" *)
  wire _00710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4618" *)
  wire _00711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4629" *)
  wire _00712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4646" *)
  wire _00713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4657" *)
  wire _00714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4674" *)
  wire _00715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9813" *)
  wire _00716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9831" *)
  wire _00717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9849" *)
  wire _00718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9867" *)
  wire _00719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4560" *)
  wire _00720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4561" *)
  wire _00721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4562" *)
  wire _00722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4563" *)
  wire _00723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4591" *)
  wire _00724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4619" *)
  wire _00725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4647" *)
  wire _00726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4675" *)
  wire _00727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4676" *)
  wire _00728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4677" *)
  wire _00729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4678" *)
  wire _00730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4679" *)
  wire _00731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4686" *)
  wire _00732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4687" *)
  wire _00733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4690" *)
  wire _00734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4691" *)
  wire _00735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4694" *)
  wire _00736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4695" *)
  wire _00737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4698" *)
  wire _00738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4699" *)
  wire _00739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4764" *)
  wire _00740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4765" *)
  wire _00741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4766" *)
  wire _00742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4767" *)
  wire _00743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4768" *)
  wire _00744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4769" *)
  wire _00745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4770" *)
  wire _00746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4771" *)
  wire _00747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4875" *)
  wire _00748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4895" *)
  wire _00749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4913" *)
  wire _00750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4931" *)
  wire _00751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4345" *)
  wire _00752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4345" *)
  wire _00753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4346" *)
  wire _00754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4347" *)
  wire _00755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4348" *)
  wire _00756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4350" *)
  wire _00757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4352" *)
  wire _00758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4356" *)
  wire _00759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4360" *)
  wire _00760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4363" *)
  wire _00761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4366" *)
  wire _00762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4369" *)
  wire _00763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4371" *)
  wire _00764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4372" *)
  wire _00765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4373" *)
  wire _00766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4398" *)
  wire _00767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4412" *)
  wire _00768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4413" *)
  wire _00769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4414" *)
  wire _00770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4417" *)
  wire _00771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4431" *)
  wire _00772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4432" *)
  wire _00773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4433" *)
  wire _00774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4436" *)
  wire _00775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4450" *)
  wire _00776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4451" *)
  wire _00777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4452" *)
  wire _00778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4455" *)
  wire _00779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4461" *)
  wire _00780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4470" *)
  wire _00781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4471" *)
  wire _00782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4474" *)
  wire _00783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4475" *)
  wire _00784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4475" *)
  wire _00785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4476" *)
  wire _00786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4481" *)
  wire _00787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4485" *)
  wire _00788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4489" *)
  wire _00789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4493" *)
  wire _00790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4495" *)
  wire _00791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4497" *)
  wire _00792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4498" *)
  wire _00793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4500" *)
  wire _00794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4501" *)
  wire _00795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4502" *)
  wire _00796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4504" *)
  wire _00797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4505" *)
  wire _00798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4506" *)
  wire _00799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4508" *)
  wire _00800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4509" *)
  wire _00801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4510" *)
  wire _00802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4512" *)
  wire _00803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4513" *)
  wire _00804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4515" *)
  wire _00805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4517" *)
  wire _00806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4519" *)
  wire _00807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4521" *)
  wire _00808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4523" *)
  wire _00809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4525" *)
  wire _00810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4527" *)
  wire _00811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4545" *)
  wire _00812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4546" *)
  wire _00813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4548" *)
  wire _00814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4550" *)
  wire _00815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *)
  wire _00816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *)
  wire _00817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *)
  wire _00818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *)
  wire _00819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *)
  wire _00820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *)
  wire _00821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *)
  wire _00822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *)
  wire _00823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4589" *)
  wire _00824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4617" *)
  wire _00825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4645" *)
  wire _00826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4673" *)
  wire _00827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4680" *)
  wire _00828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4701" *)
  wire _00829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4704" *)
  wire _00830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4705" *)
  wire _00831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4717" *)
  wire _00832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4720" *)
  wire _00833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4721" *)
  wire _00834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4733" *)
  wire _00835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4736" *)
  wire _00836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4737" *)
  wire _00837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4749" *)
  wire _00838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4752" *)
  wire _00839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4753" *)
  wire _00840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4764" *)
  wire _00841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4766" *)
  wire _00842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4768" *)
  wire _00843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4770" *)
  wire _00844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4875" *)
  wire _00845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4891" *)
  wire _00846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4895" *)
  wire _00847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4909" *)
  wire _00848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4913" *)
  wire _00849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4927" *)
  wire _00850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4931" *)
  wire _00851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4980" *)
  wire _00852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4981" *)
  wire _00853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5498" *)
  wire _00854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6014" *)
  wire _00855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6530" *)
  wire _00856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7046" *)
  wire _00857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7088" *)
  wire _00858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7091" *)
  wire _00859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7094" *)
  wire _00860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7097" *)
  wire _00861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7112" *)
  wire _00862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7127" *)
  wire _00863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7142" *)
  wire _00864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7156" *)
  wire _00865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7158" *)
  wire _00866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7296" *)
  wire _00867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7304" *)
  wire _00868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7307" *)
  wire _00869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7318" *)
  wire _00870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7319" *)
  wire _00871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7325" *)
  wire _00872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7329" *)
  wire _00873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7333" *)
  wire _00874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7342" *)
  wire _00875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7370" *)
  wire _00876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7387" *)
  wire _00877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7474" *)
  wire _00878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7482" *)
  wire _00879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7490" *)
  wire _00880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7553" *)
  wire _00881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7605" *)
  wire _00882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7657" *)
  wire _00883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7709" *)
  wire _00884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7747" *)
  wire _00885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7866" *)
  wire _00886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8003" *)
  wire _00887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8140" *)
  wire _00888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8267" *)
  wire _00889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8277" *)
  wire _00890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8383" *)
  wire _00891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8430" *)
  wire _00892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8439" *)
  wire _00893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8539" *)
  wire _00894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8605" *)
  wire _00895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8670" *)
  wire _00896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8735" *)
  wire _00897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8768" *)
  wire _00898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8776" *)
  wire _00899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8804" *)
  wire _00900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8832" *)
  wire _00901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8860" *)
  wire _00902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8880" *)
  wire _00903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8902" *)
  wire _00904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8911" *)
  wire _00905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8932" *)
  wire _00906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8954" *)
  wire _00907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8975" *)
  wire _00908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8975" *)
  wire _00909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8983" *)
  wire _00910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8991" *)
  wire _00911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8991" *)
  wire _00912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8999" *)
  wire _00913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9007" *)
  wire _00914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9007" *)
  wire _00915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9015" *)
  wire _00916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9023" *)
  wire _00917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9023" *)
  wire _00918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9031" *)
  wire _00919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9079" *)
  wire _00920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *)
  wire _00921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9098" *)
  wire _00922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *)
  wire _00923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9117" *)
  wire _00924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *)
  wire _00925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9136" *)
  wire _00926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9146" *)
  wire _00927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9155" *)
  wire _00928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9161" *)
  wire _00929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9169" *)
  wire _00930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9176" *)
  wire _00931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9184" *)
  wire _00932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9191" *)
  wire _00933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9199" *)
  wire _00934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9205" *)
  wire _00935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9213" *)
  wire _00936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9233" *)
  wire _00937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9251" *)
  wire _00938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9269" *)
  wire _00939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9287" *)
  wire _00940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9323" *)
  wire _00941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9327" *)
  wire _00942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9331" *)
  wire _00943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9338" *)
  wire _00944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9340" *)
  wire _00945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9343" *)
  wire _00946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9351" *)
  wire _00947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9357" *)
  wire _00948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9375" *)
  wire _00949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9380" *)
  wire _00950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9394" *)
  wire _00951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *)
  wire _00952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *)
  wire _00953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *)
  wire _00954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9426" *)
  wire _00955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9431" *)
  wire _00956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9435" *)
  wire _00957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9441" *)
  wire _00958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9444" *)
  wire _00959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9455" *)
  wire _00960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9461" *)
  wire _00961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9476" *)
  wire _00962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9498" *)
  wire _00963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9504" *)
  wire _00964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9507" *)
  wire _00965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9507" *)
  wire _00966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9508" *)
  wire _00967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9531" *)
  wire _00968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9536" *)
  wire _00969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9540" *)
  wire _00970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9546" *)
  wire _00971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9549" *)
  wire _00972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9560" *)
  wire _00973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9566" *)
  wire _00974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9581" *)
  wire _00975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9603" *)
  wire _00976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9609" *)
  wire _00977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9612" *)
  wire _00978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9612" *)
  wire _00979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9613" *)
  wire _00980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9636" *)
  wire _00981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9641" *)
  wire _00982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9645" *)
  wire _00983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9651" *)
  wire _00984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9654" *)
  wire _00985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9665" *)
  wire _00986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9671" *)
  wire _00987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9686" *)
  wire _00988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9709" *)
  wire _00989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9715" *)
  wire _00990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9718" *)
  wire _00991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9718" *)
  wire _00992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9719" *)
  wire _00993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9801" *)
  wire _00994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9883" *)
  wire _00995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9892" *)
  wire _00996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9901" *)
  wire _00997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9912" *)
  wire _00998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _00999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _01000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _01001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _01002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _01003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _01004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _01005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *)
  wire [7:0] _01006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _01007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _01008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _01009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _01010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _01011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _01012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _01013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *)
  wire [7:0] _01014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _01015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _01016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _01017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _01018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _01019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _01020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _01021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *)
  wire [7:0] _01022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4344" *)
  wire _01023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4345" *)
  wire _01024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4373" *)
  wire _01025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4373" *)
  wire _01026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4375" *)
  wire _01027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4375" *)
  wire _01028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4379" *)
  wire _01029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4379" *)
  wire _01030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4381" *)
  wire _01031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4381" *)
  wire _01032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4385" *)
  wire _01033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4385" *)
  wire _01034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4387" *)
  wire _01035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4387" *)
  wire _01036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4391" *)
  wire _01037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4391" *)
  wire _01038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4393" *)
  wire _01039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4393" *)
  wire _01040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4399" *)
  wire _01041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4399" *)
  wire _01042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4401" *)
  wire _01043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4401" *)
  wire _01044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4413" *)
  wire _01045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4418" *)
  wire _01046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4420" *)
  wire _01047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4422" *)
  wire _01048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4422" *)
  wire _01049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4432" *)
  wire _01050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4437" *)
  wire _01051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4439" *)
  wire _01052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4441" *)
  wire _01053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4441" *)
  wire _01054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4451" *)
  wire _01055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4456" *)
  wire _01056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4456" *)
  wire _01057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4458" *)
  wire _01058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4460" *)
  wire _01059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4460" *)
  wire _01060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4470" *)
  wire _01061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4475" *)
  wire _01062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4500" *)
  wire _01063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4500" *)
  wire _01064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4504" *)
  wire _01065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4508" *)
  wire _01066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4512" *)
  wire _01067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4531" *)
  wire _01068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4535" *)
  wire _01069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4539" *)
  wire _01070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4542" *)
  wire _01071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4544" *)
  wire _01072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *)
  wire _01073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *)
  wire _01074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *)
  wire _01075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *)
  wire _01076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *)
  wire _01077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *)
  wire _01078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *)
  wire _01079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *)
  wire _01080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *)
  wire _01081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *)
  wire _01082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *)
  wire _01083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *)
  wire _01084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4576" *)
  wire _01085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4577" *)
  wire _01086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4577" *)
  wire _01087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4578" *)
  wire _01088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4578" *)
  wire _01089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4579" *)
  wire _01090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4579" *)
  wire _01091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4580" *)
  wire _01092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4580" *)
  wire _01093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4581" *)
  wire _01094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4581" *)
  wire _01095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4582" *)
  wire _01096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4582" *)
  wire _01097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4583" *)
  wire _01098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4583" *)
  wire _01099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4584" *)
  wire _01100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4584" *)
  wire _01101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4585" *)
  wire _01102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4585" *)
  wire _01103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4586" *)
  wire _01104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4586" *)
  wire _01105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4587" *)
  wire _01106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4587" *)
  wire _01107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4589" *)
  wire _01108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4604" *)
  wire _01109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4605" *)
  wire _01110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4605" *)
  wire _01111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4606" *)
  wire _01112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4606" *)
  wire _01113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4607" *)
  wire _01114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4607" *)
  wire _01115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4608" *)
  wire _01116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4608" *)
  wire _01117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4609" *)
  wire _01118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4609" *)
  wire _01119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4610" *)
  wire _01120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4610" *)
  wire _01121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4611" *)
  wire _01122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4611" *)
  wire _01123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4612" *)
  wire _01124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4612" *)
  wire _01125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4613" *)
  wire _01126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4613" *)
  wire _01127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4614" *)
  wire _01128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4614" *)
  wire _01129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4615" *)
  wire _01130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4615" *)
  wire _01131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4617" *)
  wire _01132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4632" *)
  wire _01133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4633" *)
  wire _01134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4633" *)
  wire _01135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4634" *)
  wire _01136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4634" *)
  wire _01137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4635" *)
  wire _01138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4635" *)
  wire _01139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4636" *)
  wire _01140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4636" *)
  wire _01141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4637" *)
  wire _01142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4637" *)
  wire _01143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4638" *)
  wire _01144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4638" *)
  wire _01145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4639" *)
  wire _01146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4639" *)
  wire _01147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4640" *)
  wire _01148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4640" *)
  wire _01149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4641" *)
  wire _01150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4641" *)
  wire _01151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4642" *)
  wire _01152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4642" *)
  wire _01153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4643" *)
  wire _01154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4643" *)
  wire _01155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4645" *)
  wire _01156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4660" *)
  wire _01157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4661" *)
  wire _01158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4661" *)
  wire _01159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4662" *)
  wire _01160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4662" *)
  wire _01161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4663" *)
  wire _01162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4663" *)
  wire _01163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4664" *)
  wire _01164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4664" *)
  wire _01165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4665" *)
  wire _01166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4665" *)
  wire _01167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4666" *)
  wire _01168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4666" *)
  wire _01169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4667" *)
  wire _01170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4667" *)
  wire _01171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4668" *)
  wire _01172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4668" *)
  wire _01173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4669" *)
  wire _01174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4669" *)
  wire _01175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4670" *)
  wire _01176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4670" *)
  wire _01177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4671" *)
  wire _01178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4671" *)
  wire _01179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4673" *)
  wire _01180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4680" *)
  wire _01181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4681" *)
  wire _01182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4682" *)
  wire _01183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4683" *)
  wire _01184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4697" *)
  wire _01185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4765" *)
  wire _01186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4767" *)
  wire _01187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4769" *)
  wire _01188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4771" *)
  wire _01189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4783" *)
  wire _01190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4789" *)
  wire _01191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4804" *)
  wire _01192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4810" *)
  wire _01193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4824" *)
  wire _01194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4830" *)
  wire _01195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4844" *)
  wire _01196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4850" *)
  wire _01197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4853" *)
  wire _01198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4854" *)
  wire _01199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4855" *)
  wire _01200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4856" *)
  wire _01201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4867" *)
  wire _01202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4988" *)
  wire _01203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4988" *)
  wire _01204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4989" *)
  wire _01205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4989" *)
  wire _01206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4990" *)
  wire _01207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4990" *)
  wire _01208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4991" *)
  wire _01209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4991" *)
  wire _01210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4992" *)
  wire _01211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4992" *)
  wire _01212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4993" *)
  wire _01213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4993" *)
  wire _01214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4994" *)
  wire _01215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4994" *)
  wire _01216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4995" *)
  wire _01217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4995" *)
  wire _01218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4996" *)
  wire _01219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4996" *)
  wire _01220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4997" *)
  wire _01221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4997" *)
  wire _01222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4998" *)
  wire _01223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4998" *)
  wire _01224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4999" *)
  wire _01225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4999" *)
  wire _01226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5000" *)
  wire _01227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5000" *)
  wire _01228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5001" *)
  wire _01229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5001" *)
  wire _01230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5002" *)
  wire _01231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5002" *)
  wire _01232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5003" *)
  wire _01233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5003" *)
  wire _01234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5004" *)
  wire _01235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5004" *)
  wire _01236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5005" *)
  wire _01237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5005" *)
  wire _01238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5006" *)
  wire _01239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5006" *)
  wire _01240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5007" *)
  wire _01241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5007" *)
  wire _01242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5008" *)
  wire _01243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5008" *)
  wire _01244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5009" *)
  wire _01245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5009" *)
  wire _01246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5010" *)
  wire _01247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5010" *)
  wire _01248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5011" *)
  wire _01249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5011" *)
  wire _01250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5012" *)
  wire _01251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5012" *)
  wire _01252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5013" *)
  wire _01253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5013" *)
  wire _01254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5014" *)
  wire _01255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5014" *)
  wire _01256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5015" *)
  wire _01257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5015" *)
  wire _01258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5016" *)
  wire _01259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5016" *)
  wire _01260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5017" *)
  wire _01261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5017" *)
  wire _01262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5018" *)
  wire _01263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5018" *)
  wire _01264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5019" *)
  wire _01265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5019" *)
  wire _01266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5020" *)
  wire _01267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5020" *)
  wire _01268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5021" *)
  wire _01269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5021" *)
  wire _01270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5022" *)
  wire _01271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5022" *)
  wire _01272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5023" *)
  wire _01273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5023" *)
  wire _01274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5024" *)
  wire _01275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5024" *)
  wire _01276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5025" *)
  wire _01277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5025" *)
  wire _01278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5026" *)
  wire _01279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5026" *)
  wire _01280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5027" *)
  wire _01281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5027" *)
  wire _01282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5028" *)
  wire _01283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5028" *)
  wire _01284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5029" *)
  wire _01285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5029" *)
  wire _01286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5030" *)
  wire _01287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5030" *)
  wire _01288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5031" *)
  wire _01289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5031" *)
  wire _01290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5032" *)
  wire _01291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5032" *)
  wire _01292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5033" *)
  wire _01293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5033" *)
  wire _01294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5034" *)
  wire _01295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5034" *)
  wire _01296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5035" *)
  wire _01297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5035" *)
  wire _01298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5036" *)
  wire _01299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5036" *)
  wire _01300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5037" *)
  wire _01301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5037" *)
  wire _01302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5038" *)
  wire _01303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5038" *)
  wire _01304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5039" *)
  wire _01305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5039" *)
  wire _01306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5040" *)
  wire _01307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5040" *)
  wire _01308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5041" *)
  wire _01309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5041" *)
  wire _01310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5042" *)
  wire _01311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5042" *)
  wire _01312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5043" *)
  wire _01313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5043" *)
  wire _01314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5044" *)
  wire _01315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5044" *)
  wire _01316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5045" *)
  wire _01317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5045" *)
  wire _01318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5046" *)
  wire _01319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5046" *)
  wire _01320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5047" *)
  wire _01321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5047" *)
  wire _01322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5048" *)
  wire _01323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5048" *)
  wire _01324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5049" *)
  wire _01325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5049" *)
  wire _01326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5050" *)
  wire _01327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5050" *)
  wire _01328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5051" *)
  wire _01329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5051" *)
  wire _01330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5052" *)
  wire _01331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5052" *)
  wire _01332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5053" *)
  wire _01333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5053" *)
  wire _01334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5054" *)
  wire _01335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5054" *)
  wire _01336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5055" *)
  wire _01337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5055" *)
  wire _01338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5056" *)
  wire _01339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5056" *)
  wire _01340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5057" *)
  wire _01341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5057" *)
  wire _01342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5058" *)
  wire _01343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5058" *)
  wire _01344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5059" *)
  wire _01345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5059" *)
  wire _01346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5060" *)
  wire _01347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5060" *)
  wire _01348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5061" *)
  wire _01349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5061" *)
  wire _01350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5062" *)
  wire _01351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5062" *)
  wire _01352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5063" *)
  wire _01353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5063" *)
  wire _01354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5064" *)
  wire _01355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5064" *)
  wire _01356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5065" *)
  wire _01357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5065" *)
  wire _01358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5066" *)
  wire _01359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5066" *)
  wire _01360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5067" *)
  wire _01361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5067" *)
  wire _01362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5068" *)
  wire _01363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5068" *)
  wire _01364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5069" *)
  wire _01365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5069" *)
  wire _01366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5070" *)
  wire _01367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5070" *)
  wire _01368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5071" *)
  wire _01369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5071" *)
  wire _01370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5072" *)
  wire _01371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5072" *)
  wire _01372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5073" *)
  wire _01373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5073" *)
  wire _01374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5074" *)
  wire _01375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5074" *)
  wire _01376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5075" *)
  wire _01377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5075" *)
  wire _01378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5076" *)
  wire _01379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5076" *)
  wire _01380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5077" *)
  wire _01381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5077" *)
  wire _01382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5078" *)
  wire _01383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5078" *)
  wire _01384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5079" *)
  wire _01385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5079" *)
  wire _01386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5080" *)
  wire _01387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5080" *)
  wire _01388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5081" *)
  wire _01389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5081" *)
  wire _01390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5082" *)
  wire _01391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5082" *)
  wire _01392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5083" *)
  wire _01393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5083" *)
  wire _01394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5084" *)
  wire _01395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5084" *)
  wire _01396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5085" *)
  wire _01397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5085" *)
  wire _01398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5086" *)
  wire _01399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5086" *)
  wire _01400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5087" *)
  wire _01401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5087" *)
  wire _01402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5088" *)
  wire _01403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5088" *)
  wire _01404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5089" *)
  wire _01405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5089" *)
  wire _01406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5090" *)
  wire _01407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5090" *)
  wire _01408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5091" *)
  wire _01409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5091" *)
  wire _01410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5092" *)
  wire _01411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5092" *)
  wire _01412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5093" *)
  wire _01413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5093" *)
  wire _01414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5094" *)
  wire _01415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5094" *)
  wire _01416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5095" *)
  wire _01417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5095" *)
  wire _01418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5096" *)
  wire _01419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5096" *)
  wire _01420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5097" *)
  wire _01421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5097" *)
  wire _01422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5098" *)
  wire _01423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5098" *)
  wire _01424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5099" *)
  wire _01425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5099" *)
  wire _01426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5100" *)
  wire _01427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5100" *)
  wire _01428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5101" *)
  wire _01429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5101" *)
  wire _01430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5102" *)
  wire _01431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5102" *)
  wire _01432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5103" *)
  wire _01433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5103" *)
  wire _01434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5104" *)
  wire _01435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5104" *)
  wire _01436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5105" *)
  wire _01437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5105" *)
  wire _01438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5106" *)
  wire _01439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5106" *)
  wire _01440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5107" *)
  wire _01441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5107" *)
  wire _01442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5108" *)
  wire _01443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5108" *)
  wire _01444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5109" *)
  wire _01445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5109" *)
  wire _01446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5110" *)
  wire _01447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5110" *)
  wire _01448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5111" *)
  wire _01449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5111" *)
  wire _01450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5112" *)
  wire _01451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5112" *)
  wire _01452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5113" *)
  wire _01453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5113" *)
  wire _01454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5114" *)
  wire _01455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5114" *)
  wire _01456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5115" *)
  wire _01457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5115" *)
  wire _01458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5116" *)
  wire _01459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5116" *)
  wire _01460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5117" *)
  wire _01461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5117" *)
  wire _01462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5118" *)
  wire _01463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5118" *)
  wire _01464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5119" *)
  wire _01465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5119" *)
  wire _01466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5120" *)
  wire _01467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5120" *)
  wire _01468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5121" *)
  wire _01469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5121" *)
  wire _01470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5122" *)
  wire _01471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5122" *)
  wire _01472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5123" *)
  wire _01473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5123" *)
  wire _01474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5124" *)
  wire _01475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5124" *)
  wire _01476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5125" *)
  wire _01477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5125" *)
  wire _01478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5126" *)
  wire _01479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5126" *)
  wire _01480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5127" *)
  wire _01481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5127" *)
  wire _01482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5128" *)
  wire _01483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5128" *)
  wire _01484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5129" *)
  wire _01485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5129" *)
  wire _01486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5130" *)
  wire _01487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5130" *)
  wire _01488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5131" *)
  wire _01489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5131" *)
  wire _01490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5132" *)
  wire _01491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5132" *)
  wire _01492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5133" *)
  wire _01493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5133" *)
  wire _01494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5134" *)
  wire _01495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5134" *)
  wire _01496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5135" *)
  wire _01497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5135" *)
  wire _01498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5136" *)
  wire _01499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5136" *)
  wire _01500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5137" *)
  wire _01501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5137" *)
  wire _01502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5138" *)
  wire _01503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5138" *)
  wire _01504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5139" *)
  wire _01505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5139" *)
  wire _01506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5140" *)
  wire _01507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5140" *)
  wire _01508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5141" *)
  wire _01509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5141" *)
  wire _01510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5142" *)
  wire _01511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5142" *)
  wire _01512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5143" *)
  wire _01513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5143" *)
  wire _01514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5144" *)
  wire _01515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5144" *)
  wire _01516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5145" *)
  wire _01517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5145" *)
  wire _01518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5146" *)
  wire _01519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5146" *)
  wire _01520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5147" *)
  wire _01521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5147" *)
  wire _01522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5148" *)
  wire _01523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5148" *)
  wire _01524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5149" *)
  wire _01525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5149" *)
  wire _01526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5150" *)
  wire _01527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5150" *)
  wire _01528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5151" *)
  wire _01529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5151" *)
  wire _01530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5152" *)
  wire _01531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5152" *)
  wire _01532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5153" *)
  wire _01533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5153" *)
  wire _01534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5154" *)
  wire _01535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5154" *)
  wire _01536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5155" *)
  wire _01537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5155" *)
  wire _01538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5156" *)
  wire _01539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5156" *)
  wire _01540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5157" *)
  wire _01541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5157" *)
  wire _01542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5158" *)
  wire _01543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5158" *)
  wire _01544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5159" *)
  wire _01545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5159" *)
  wire _01546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5160" *)
  wire _01547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5160" *)
  wire _01548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5161" *)
  wire _01549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5161" *)
  wire _01550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5162" *)
  wire _01551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5162" *)
  wire _01552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5163" *)
  wire _01553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5163" *)
  wire _01554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5164" *)
  wire _01555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5164" *)
  wire _01556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5165" *)
  wire _01557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5165" *)
  wire _01558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5166" *)
  wire _01559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5166" *)
  wire _01560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5167" *)
  wire _01561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5167" *)
  wire _01562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5168" *)
  wire _01563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5168" *)
  wire _01564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5169" *)
  wire _01565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5169" *)
  wire _01566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5170" *)
  wire _01567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5170" *)
  wire _01568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5171" *)
  wire _01569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5171" *)
  wire _01570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5172" *)
  wire _01571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5172" *)
  wire _01572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5173" *)
  wire _01573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5173" *)
  wire _01574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5174" *)
  wire _01575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5174" *)
  wire _01576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5175" *)
  wire _01577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5175" *)
  wire _01578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5176" *)
  wire _01579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5176" *)
  wire _01580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5177" *)
  wire _01581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5177" *)
  wire _01582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5178" *)
  wire _01583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5178" *)
  wire _01584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5179" *)
  wire _01585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5179" *)
  wire _01586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5180" *)
  wire _01587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5180" *)
  wire _01588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5181" *)
  wire _01589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5181" *)
  wire _01590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5182" *)
  wire _01591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5182" *)
  wire _01592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5183" *)
  wire _01593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5183" *)
  wire _01594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5184" *)
  wire _01595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5184" *)
  wire _01596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5185" *)
  wire _01597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5185" *)
  wire _01598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5186" *)
  wire _01599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5186" *)
  wire _01600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5187" *)
  wire _01601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5187" *)
  wire _01602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5188" *)
  wire _01603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5188" *)
  wire _01604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5189" *)
  wire _01605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5189" *)
  wire _01606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5190" *)
  wire _01607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5190" *)
  wire _01608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5191" *)
  wire _01609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5191" *)
  wire _01610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5192" *)
  wire _01611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5192" *)
  wire _01612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5193" *)
  wire _01613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5193" *)
  wire _01614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5194" *)
  wire _01615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5194" *)
  wire _01616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5195" *)
  wire _01617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5195" *)
  wire _01618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5196" *)
  wire _01619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5196" *)
  wire _01620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5197" *)
  wire _01621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5197" *)
  wire _01622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5198" *)
  wire _01623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5198" *)
  wire _01624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5199" *)
  wire _01625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5199" *)
  wire _01626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5200" *)
  wire _01627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5200" *)
  wire _01628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5201" *)
  wire _01629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5201" *)
  wire _01630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5202" *)
  wire _01631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5202" *)
  wire _01632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5203" *)
  wire _01633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5203" *)
  wire _01634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5204" *)
  wire _01635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5204" *)
  wire _01636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5205" *)
  wire _01637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5205" *)
  wire _01638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5206" *)
  wire _01639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5206" *)
  wire _01640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5207" *)
  wire _01641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5207" *)
  wire _01642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5208" *)
  wire _01643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5208" *)
  wire _01644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5209" *)
  wire _01645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5209" *)
  wire _01646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5210" *)
  wire _01647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5210" *)
  wire _01648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5211" *)
  wire _01649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5211" *)
  wire _01650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5212" *)
  wire _01651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5212" *)
  wire _01652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5213" *)
  wire _01653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5213" *)
  wire _01654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5214" *)
  wire _01655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5214" *)
  wire _01656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5215" *)
  wire _01657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5215" *)
  wire _01658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5216" *)
  wire _01659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5216" *)
  wire _01660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5217" *)
  wire _01661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5217" *)
  wire _01662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5218" *)
  wire _01663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5218" *)
  wire _01664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5219" *)
  wire _01665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5219" *)
  wire _01666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5220" *)
  wire _01667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5220" *)
  wire _01668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5221" *)
  wire _01669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5221" *)
  wire _01670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5222" *)
  wire _01671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5222" *)
  wire _01672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5223" *)
  wire _01673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5223" *)
  wire _01674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5224" *)
  wire _01675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5224" *)
  wire _01676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5225" *)
  wire _01677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5225" *)
  wire _01678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5226" *)
  wire _01679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5226" *)
  wire _01680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5227" *)
  wire _01681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5227" *)
  wire _01682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5228" *)
  wire _01683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5228" *)
  wire _01684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5229" *)
  wire _01685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5229" *)
  wire _01686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5230" *)
  wire _01687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5230" *)
  wire _01688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5231" *)
  wire _01689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5231" *)
  wire _01690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5232" *)
  wire _01691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5232" *)
  wire _01692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5233" *)
  wire _01693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5233" *)
  wire _01694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5234" *)
  wire _01695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5234" *)
  wire _01696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5235" *)
  wire _01697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5235" *)
  wire _01698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5236" *)
  wire _01699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5236" *)
  wire _01700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5237" *)
  wire _01701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5237" *)
  wire _01702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5238" *)
  wire _01703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5238" *)
  wire _01704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5239" *)
  wire _01705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5239" *)
  wire _01706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5240" *)
  wire _01707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5240" *)
  wire _01708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5241" *)
  wire _01709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5241" *)
  wire _01710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5242" *)
  wire _01711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5242" *)
  wire _01712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5243" *)
  wire _01713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5243" *)
  wire _01714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5244" *)
  wire _01715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5244" *)
  wire _01716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5245" *)
  wire _01717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5245" *)
  wire _01718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5246" *)
  wire _01719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5246" *)
  wire _01720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5247" *)
  wire _01721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5247" *)
  wire _01722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5248" *)
  wire _01723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5248" *)
  wire _01724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5249" *)
  wire _01725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5249" *)
  wire _01726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5250" *)
  wire _01727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5250" *)
  wire _01728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5251" *)
  wire _01729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5251" *)
  wire _01730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5252" *)
  wire _01731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5252" *)
  wire _01732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5253" *)
  wire _01733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5253" *)
  wire _01734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5254" *)
  wire _01735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5254" *)
  wire _01736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5255" *)
  wire _01737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5255" *)
  wire _01738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5256" *)
  wire _01739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5256" *)
  wire _01740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5257" *)
  wire _01741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5257" *)
  wire _01742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5258" *)
  wire _01743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5258" *)
  wire _01744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5259" *)
  wire _01745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5259" *)
  wire _01746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5260" *)
  wire _01747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5260" *)
  wire _01748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5261" *)
  wire _01749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5261" *)
  wire _01750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5262" *)
  wire _01751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5262" *)
  wire _01752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5263" *)
  wire _01753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5263" *)
  wire _01754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5264" *)
  wire _01755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5264" *)
  wire _01756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5265" *)
  wire _01757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5265" *)
  wire _01758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5266" *)
  wire _01759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5266" *)
  wire _01760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5267" *)
  wire _01761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5267" *)
  wire _01762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5268" *)
  wire _01763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5268" *)
  wire _01764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5269" *)
  wire _01765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5269" *)
  wire _01766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5270" *)
  wire _01767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5270" *)
  wire _01768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5271" *)
  wire _01769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5271" *)
  wire _01770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5272" *)
  wire _01771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5272" *)
  wire _01772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5273" *)
  wire _01773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5273" *)
  wire _01774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5274" *)
  wire _01775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5274" *)
  wire _01776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5275" *)
  wire _01777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5275" *)
  wire _01778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5276" *)
  wire _01779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5276" *)
  wire _01780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5277" *)
  wire _01781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5277" *)
  wire _01782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5278" *)
  wire _01783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5278" *)
  wire _01784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5279" *)
  wire _01785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5279" *)
  wire _01786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5280" *)
  wire _01787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5280" *)
  wire _01788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5281" *)
  wire _01789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5281" *)
  wire _01790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5282" *)
  wire _01791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5282" *)
  wire _01792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5283" *)
  wire _01793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5283" *)
  wire _01794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5284" *)
  wire _01795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5284" *)
  wire _01796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5285" *)
  wire _01797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5285" *)
  wire _01798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5286" *)
  wire _01799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5286" *)
  wire _01800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5287" *)
  wire _01801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5287" *)
  wire _01802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5288" *)
  wire _01803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5288" *)
  wire _01804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5289" *)
  wire _01805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5289" *)
  wire _01806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5290" *)
  wire _01807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5290" *)
  wire _01808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5291" *)
  wire _01809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5291" *)
  wire _01810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5292" *)
  wire _01811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5292" *)
  wire _01812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5293" *)
  wire _01813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5293" *)
  wire _01814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5294" *)
  wire _01815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5294" *)
  wire _01816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5295" *)
  wire _01817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5295" *)
  wire _01818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5296" *)
  wire _01819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5296" *)
  wire _01820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5297" *)
  wire _01821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5297" *)
  wire _01822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5298" *)
  wire _01823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5298" *)
  wire _01824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5299" *)
  wire _01825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5299" *)
  wire _01826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5300" *)
  wire _01827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5300" *)
  wire _01828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5301" *)
  wire _01829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5301" *)
  wire _01830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5302" *)
  wire _01831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5302" *)
  wire _01832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5303" *)
  wire _01833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5303" *)
  wire _01834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5304" *)
  wire _01835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5304" *)
  wire _01836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5305" *)
  wire _01837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5305" *)
  wire _01838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5306" *)
  wire _01839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5306" *)
  wire _01840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5307" *)
  wire _01841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5307" *)
  wire _01842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5308" *)
  wire _01843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5308" *)
  wire _01844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5309" *)
  wire _01845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5309" *)
  wire _01846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5310" *)
  wire _01847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5310" *)
  wire _01848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5311" *)
  wire _01849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5311" *)
  wire _01850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5312" *)
  wire _01851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5312" *)
  wire _01852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5313" *)
  wire _01853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5313" *)
  wire _01854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5314" *)
  wire _01855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5314" *)
  wire _01856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5315" *)
  wire _01857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5315" *)
  wire _01858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5316" *)
  wire _01859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5316" *)
  wire _01860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5317" *)
  wire _01861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5317" *)
  wire _01862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5318" *)
  wire _01863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5318" *)
  wire _01864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5319" *)
  wire _01865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5319" *)
  wire _01866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5320" *)
  wire _01867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5320" *)
  wire _01868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5321" *)
  wire _01869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5321" *)
  wire _01870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5322" *)
  wire _01871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5322" *)
  wire _01872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5323" *)
  wire _01873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5323" *)
  wire _01874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5324" *)
  wire _01875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5324" *)
  wire _01876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5325" *)
  wire _01877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5325" *)
  wire _01878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5326" *)
  wire _01879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5326" *)
  wire _01880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5327" *)
  wire _01881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5327" *)
  wire _01882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5328" *)
  wire _01883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5328" *)
  wire _01884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5329" *)
  wire _01885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5329" *)
  wire _01886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5330" *)
  wire _01887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5330" *)
  wire _01888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5331" *)
  wire _01889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5331" *)
  wire _01890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5332" *)
  wire _01891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5332" *)
  wire _01892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5333" *)
  wire _01893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5333" *)
  wire _01894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5334" *)
  wire _01895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5334" *)
  wire _01896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5335" *)
  wire _01897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5335" *)
  wire _01898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5336" *)
  wire _01899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5336" *)
  wire _01900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5337" *)
  wire _01901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5337" *)
  wire _01902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5338" *)
  wire _01903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5338" *)
  wire _01904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5339" *)
  wire _01905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5339" *)
  wire _01906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5340" *)
  wire _01907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5340" *)
  wire _01908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5341" *)
  wire _01909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5341" *)
  wire _01910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5342" *)
  wire _01911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5342" *)
  wire _01912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5343" *)
  wire _01913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5343" *)
  wire _01914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5344" *)
  wire _01915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5344" *)
  wire _01916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5345" *)
  wire _01917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5345" *)
  wire _01918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5346" *)
  wire _01919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5346" *)
  wire _01920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5347" *)
  wire _01921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5347" *)
  wire _01922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5348" *)
  wire _01923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5348" *)
  wire _01924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5349" *)
  wire _01925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5349" *)
  wire _01926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5350" *)
  wire _01927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5350" *)
  wire _01928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5351" *)
  wire _01929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5351" *)
  wire _01930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5352" *)
  wire _01931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5352" *)
  wire _01932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5353" *)
  wire _01933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5353" *)
  wire _01934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5354" *)
  wire _01935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5354" *)
  wire _01936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5355" *)
  wire _01937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5355" *)
  wire _01938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5356" *)
  wire _01939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5356" *)
  wire _01940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5357" *)
  wire _01941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5357" *)
  wire _01942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5358" *)
  wire _01943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5358" *)
  wire _01944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5359" *)
  wire _01945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5359" *)
  wire _01946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5360" *)
  wire _01947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5360" *)
  wire _01948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5361" *)
  wire _01949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5361" *)
  wire _01950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5362" *)
  wire _01951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5362" *)
  wire _01952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5363" *)
  wire _01953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5363" *)
  wire _01954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5364" *)
  wire _01955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5364" *)
  wire _01956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5365" *)
  wire _01957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5365" *)
  wire _01958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5366" *)
  wire _01959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5366" *)
  wire _01960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5367" *)
  wire _01961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5367" *)
  wire _01962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5368" *)
  wire _01963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5368" *)
  wire _01964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5369" *)
  wire _01965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5369" *)
  wire _01966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5370" *)
  wire _01967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5370" *)
  wire _01968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5371" *)
  wire _01969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5371" *)
  wire _01970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5372" *)
  wire _01971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5372" *)
  wire _01972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5373" *)
  wire _01973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5373" *)
  wire _01974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5374" *)
  wire _01975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5374" *)
  wire _01976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5375" *)
  wire _01977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5375" *)
  wire _01978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5376" *)
  wire _01979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5376" *)
  wire _01980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5377" *)
  wire _01981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5377" *)
  wire _01982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5378" *)
  wire _01983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5378" *)
  wire _01984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5379" *)
  wire _01985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5379" *)
  wire _01986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5380" *)
  wire _01987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5380" *)
  wire _01988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5381" *)
  wire _01989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5381" *)
  wire _01990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5382" *)
  wire _01991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5382" *)
  wire _01992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5383" *)
  wire _01993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5383" *)
  wire _01994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5384" *)
  wire _01995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5384" *)
  wire _01996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5385" *)
  wire _01997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5385" *)
  wire _01998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5386" *)
  wire _01999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5386" *)
  wire _02000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5387" *)
  wire _02001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5387" *)
  wire _02002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5388" *)
  wire _02003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5388" *)
  wire _02004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5389" *)
  wire _02005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5389" *)
  wire _02006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5390" *)
  wire _02007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5390" *)
  wire _02008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5391" *)
  wire _02009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5391" *)
  wire _02010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5392" *)
  wire _02011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5392" *)
  wire _02012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5393" *)
  wire _02013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5393" *)
  wire _02014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5394" *)
  wire _02015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5394" *)
  wire _02016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5395" *)
  wire _02017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5395" *)
  wire _02018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5396" *)
  wire _02019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5396" *)
  wire _02020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5397" *)
  wire _02021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5397" *)
  wire _02022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5398" *)
  wire _02023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5398" *)
  wire _02024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5399" *)
  wire _02025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5399" *)
  wire _02026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5400" *)
  wire _02027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5400" *)
  wire _02028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5401" *)
  wire _02029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5401" *)
  wire _02030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5402" *)
  wire _02031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5402" *)
  wire _02032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5403" *)
  wire _02033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5403" *)
  wire _02034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5404" *)
  wire _02035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5404" *)
  wire _02036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5405" *)
  wire _02037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5405" *)
  wire _02038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5406" *)
  wire _02039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5406" *)
  wire _02040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5407" *)
  wire _02041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5407" *)
  wire _02042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5408" *)
  wire _02043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5408" *)
  wire _02044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5409" *)
  wire _02045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5409" *)
  wire _02046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5410" *)
  wire _02047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5410" *)
  wire _02048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5411" *)
  wire _02049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5411" *)
  wire _02050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5412" *)
  wire _02051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5412" *)
  wire _02052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5413" *)
  wire _02053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5413" *)
  wire _02054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5414" *)
  wire _02055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5414" *)
  wire _02056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5415" *)
  wire _02057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5415" *)
  wire _02058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5416" *)
  wire _02059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5416" *)
  wire _02060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5417" *)
  wire _02061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5417" *)
  wire _02062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5418" *)
  wire _02063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5418" *)
  wire _02064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5419" *)
  wire _02065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5419" *)
  wire _02066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5420" *)
  wire _02067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5420" *)
  wire _02068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5421" *)
  wire _02069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5421" *)
  wire _02070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5422" *)
  wire _02071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5422" *)
  wire _02072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5423" *)
  wire _02073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5423" *)
  wire _02074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5424" *)
  wire _02075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5424" *)
  wire _02076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5425" *)
  wire _02077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5425" *)
  wire _02078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5426" *)
  wire _02079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5426" *)
  wire _02080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5427" *)
  wire _02081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5427" *)
  wire _02082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5428" *)
  wire _02083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5428" *)
  wire _02084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5429" *)
  wire _02085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5429" *)
  wire _02086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5430" *)
  wire _02087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5430" *)
  wire _02088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5431" *)
  wire _02089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5431" *)
  wire _02090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5432" *)
  wire _02091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5432" *)
  wire _02092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5433" *)
  wire _02093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5433" *)
  wire _02094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5434" *)
  wire _02095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5434" *)
  wire _02096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5435" *)
  wire _02097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5435" *)
  wire _02098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5436" *)
  wire _02099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5436" *)
  wire _02100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5437" *)
  wire _02101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5437" *)
  wire _02102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5438" *)
  wire _02103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5438" *)
  wire _02104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5439" *)
  wire _02105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5439" *)
  wire _02106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5440" *)
  wire _02107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5440" *)
  wire _02108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5441" *)
  wire _02109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5441" *)
  wire _02110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5442" *)
  wire _02111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5442" *)
  wire _02112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5443" *)
  wire _02113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5443" *)
  wire _02114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5444" *)
  wire _02115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5444" *)
  wire _02116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5445" *)
  wire _02117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5445" *)
  wire _02118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5446" *)
  wire _02119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5446" *)
  wire _02120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5447" *)
  wire _02121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5447" *)
  wire _02122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5448" *)
  wire _02123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5448" *)
  wire _02124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5449" *)
  wire _02125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5449" *)
  wire _02126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5450" *)
  wire _02127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5450" *)
  wire _02128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5451" *)
  wire _02129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5451" *)
  wire _02130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5452" *)
  wire _02131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5452" *)
  wire _02132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5453" *)
  wire _02133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5453" *)
  wire _02134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5454" *)
  wire _02135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5454" *)
  wire _02136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5455" *)
  wire _02137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5455" *)
  wire _02138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5456" *)
  wire _02139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5456" *)
  wire _02140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5457" *)
  wire _02141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5457" *)
  wire _02142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5458" *)
  wire _02143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5458" *)
  wire _02144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5459" *)
  wire _02145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5459" *)
  wire _02146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5460" *)
  wire _02147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5460" *)
  wire _02148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5461" *)
  wire _02149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5461" *)
  wire _02150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5462" *)
  wire _02151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5462" *)
  wire _02152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5463" *)
  wire _02153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5463" *)
  wire _02154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5464" *)
  wire _02155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5464" *)
  wire _02156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5465" *)
  wire _02157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5465" *)
  wire _02158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5466" *)
  wire _02159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5466" *)
  wire _02160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5467" *)
  wire _02161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5467" *)
  wire _02162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5468" *)
  wire _02163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5468" *)
  wire _02164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5469" *)
  wire _02165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5469" *)
  wire _02166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5470" *)
  wire _02167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5470" *)
  wire _02168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5471" *)
  wire _02169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5471" *)
  wire _02170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5472" *)
  wire _02171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5472" *)
  wire _02172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5473" *)
  wire _02173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5473" *)
  wire _02174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5474" *)
  wire _02175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5474" *)
  wire _02176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5475" *)
  wire _02177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5475" *)
  wire _02178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5476" *)
  wire _02179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5476" *)
  wire _02180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5477" *)
  wire _02181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5477" *)
  wire _02182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5478" *)
  wire _02183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5478" *)
  wire _02184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5479" *)
  wire _02185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5479" *)
  wire _02186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5480" *)
  wire _02187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5480" *)
  wire _02188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5481" *)
  wire _02189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5481" *)
  wire _02190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5482" *)
  wire _02191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5482" *)
  wire _02192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5483" *)
  wire _02193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5483" *)
  wire _02194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5484" *)
  wire _02195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5484" *)
  wire _02196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5485" *)
  wire _02197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5485" *)
  wire _02198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5486" *)
  wire _02199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5486" *)
  wire _02200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5487" *)
  wire _02201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5487" *)
  wire _02202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5488" *)
  wire _02203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5488" *)
  wire _02204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5489" *)
  wire _02205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5489" *)
  wire _02206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5490" *)
  wire _02207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5490" *)
  wire _02208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5491" *)
  wire _02209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5491" *)
  wire _02210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5492" *)
  wire _02211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5492" *)
  wire _02212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5493" *)
  wire _02213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5493" *)
  wire _02214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5494" *)
  wire _02215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5494" *)
  wire _02216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5495" *)
  wire _02217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5495" *)
  wire _02218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5496" *)
  wire _02219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5496" *)
  wire _02220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5497" *)
  wire _02221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5497" *)
  wire _02222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5498" *)
  wire _02223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5498" *)
  wire _02224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5504" *)
  wire _02225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5504" *)
  wire _02226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5505" *)
  wire _02227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5505" *)
  wire _02228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5506" *)
  wire _02229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5506" *)
  wire _02230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5507" *)
  wire _02231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5507" *)
  wire _02232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5508" *)
  wire _02233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5508" *)
  wire _02234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5509" *)
  wire _02235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5509" *)
  wire _02236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5510" *)
  wire _02237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5510" *)
  wire _02238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5511" *)
  wire _02239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5511" *)
  wire _02240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5512" *)
  wire _02241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5512" *)
  wire _02242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5513" *)
  wire _02243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5513" *)
  wire _02244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5514" *)
  wire _02245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5514" *)
  wire _02246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5515" *)
  wire _02247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5515" *)
  wire _02248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5516" *)
  wire _02249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5516" *)
  wire _02250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5517" *)
  wire _02251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5517" *)
  wire _02252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5518" *)
  wire _02253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5518" *)
  wire _02254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5519" *)
  wire _02255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5519" *)
  wire _02256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5520" *)
  wire _02257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5520" *)
  wire _02258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5521" *)
  wire _02259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5521" *)
  wire _02260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5522" *)
  wire _02261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5522" *)
  wire _02262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5523" *)
  wire _02263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5523" *)
  wire _02264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5524" *)
  wire _02265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5524" *)
  wire _02266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5525" *)
  wire _02267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5525" *)
  wire _02268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5526" *)
  wire _02269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5526" *)
  wire _02270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5527" *)
  wire _02271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5527" *)
  wire _02272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5528" *)
  wire _02273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5528" *)
  wire _02274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5529" *)
  wire _02275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5529" *)
  wire _02276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5530" *)
  wire _02277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5530" *)
  wire _02278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5531" *)
  wire _02279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5531" *)
  wire _02280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5532" *)
  wire _02281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5532" *)
  wire _02282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5533" *)
  wire _02283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5533" *)
  wire _02284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5534" *)
  wire _02285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5534" *)
  wire _02286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5535" *)
  wire _02287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5535" *)
  wire _02288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5536" *)
  wire _02289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5536" *)
  wire _02290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5537" *)
  wire _02291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5537" *)
  wire _02292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5538" *)
  wire _02293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5538" *)
  wire _02294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5539" *)
  wire _02295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5539" *)
  wire _02296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5540" *)
  wire _02297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5540" *)
  wire _02298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5541" *)
  wire _02299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5541" *)
  wire _02300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5542" *)
  wire _02301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5542" *)
  wire _02302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5543" *)
  wire _02303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5543" *)
  wire _02304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5544" *)
  wire _02305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5544" *)
  wire _02306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5545" *)
  wire _02307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5545" *)
  wire _02308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5546" *)
  wire _02309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5546" *)
  wire _02310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5547" *)
  wire _02311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5547" *)
  wire _02312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5548" *)
  wire _02313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5548" *)
  wire _02314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5549" *)
  wire _02315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5549" *)
  wire _02316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5550" *)
  wire _02317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5550" *)
  wire _02318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5551" *)
  wire _02319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5551" *)
  wire _02320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5552" *)
  wire _02321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5552" *)
  wire _02322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5553" *)
  wire _02323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5553" *)
  wire _02324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5554" *)
  wire _02325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5554" *)
  wire _02326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5555" *)
  wire _02327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5555" *)
  wire _02328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5556" *)
  wire _02329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5556" *)
  wire _02330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5557" *)
  wire _02331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5557" *)
  wire _02332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5558" *)
  wire _02333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5558" *)
  wire _02334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5559" *)
  wire _02335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5559" *)
  wire _02336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5560" *)
  wire _02337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5560" *)
  wire _02338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5561" *)
  wire _02339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5561" *)
  wire _02340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5562" *)
  wire _02341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5562" *)
  wire _02342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5563" *)
  wire _02343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5563" *)
  wire _02344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5564" *)
  wire _02345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5564" *)
  wire _02346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5565" *)
  wire _02347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5565" *)
  wire _02348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5566" *)
  wire _02349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5566" *)
  wire _02350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5567" *)
  wire _02351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5567" *)
  wire _02352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5568" *)
  wire _02353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5568" *)
  wire _02354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5569" *)
  wire _02355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5569" *)
  wire _02356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5570" *)
  wire _02357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5570" *)
  wire _02358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5571" *)
  wire _02359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5571" *)
  wire _02360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5572" *)
  wire _02361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5572" *)
  wire _02362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5573" *)
  wire _02363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5573" *)
  wire _02364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5574" *)
  wire _02365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5574" *)
  wire _02366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5575" *)
  wire _02367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5575" *)
  wire _02368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5576" *)
  wire _02369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5576" *)
  wire _02370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5577" *)
  wire _02371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5577" *)
  wire _02372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5578" *)
  wire _02373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5578" *)
  wire _02374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5579" *)
  wire _02375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5579" *)
  wire _02376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5580" *)
  wire _02377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5580" *)
  wire _02378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5581" *)
  wire _02379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5581" *)
  wire _02380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5582" *)
  wire _02381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5582" *)
  wire _02382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5583" *)
  wire _02383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5583" *)
  wire _02384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5584" *)
  wire _02385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5584" *)
  wire _02386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5585" *)
  wire _02387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5585" *)
  wire _02388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5586" *)
  wire _02389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5586" *)
  wire _02390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5587" *)
  wire _02391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5587" *)
  wire _02392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5588" *)
  wire _02393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5588" *)
  wire _02394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5589" *)
  wire _02395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5589" *)
  wire _02396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5590" *)
  wire _02397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5590" *)
  wire _02398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5591" *)
  wire _02399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5591" *)
  wire _02400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5592" *)
  wire _02401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5592" *)
  wire _02402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5593" *)
  wire _02403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5593" *)
  wire _02404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5594" *)
  wire _02405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5594" *)
  wire _02406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5595" *)
  wire _02407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5595" *)
  wire _02408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5596" *)
  wire _02409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5596" *)
  wire _02410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5597" *)
  wire _02411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5597" *)
  wire _02412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5598" *)
  wire _02413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5598" *)
  wire _02414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5599" *)
  wire _02415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5599" *)
  wire _02416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5600" *)
  wire _02417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5600" *)
  wire _02418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5601" *)
  wire _02419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5601" *)
  wire _02420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5602" *)
  wire _02421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5602" *)
  wire _02422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5603" *)
  wire _02423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5603" *)
  wire _02424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5604" *)
  wire _02425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5604" *)
  wire _02426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5605" *)
  wire _02427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5605" *)
  wire _02428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5606" *)
  wire _02429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5606" *)
  wire _02430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5607" *)
  wire _02431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5607" *)
  wire _02432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5608" *)
  wire _02433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5608" *)
  wire _02434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5609" *)
  wire _02435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5609" *)
  wire _02436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5610" *)
  wire _02437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5610" *)
  wire _02438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5611" *)
  wire _02439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5611" *)
  wire _02440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5612" *)
  wire _02441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5612" *)
  wire _02442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5613" *)
  wire _02443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5613" *)
  wire _02444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5614" *)
  wire _02445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5614" *)
  wire _02446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5615" *)
  wire _02447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5615" *)
  wire _02448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5616" *)
  wire _02449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5616" *)
  wire _02450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5617" *)
  wire _02451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5617" *)
  wire _02452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5618" *)
  wire _02453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5618" *)
  wire _02454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5619" *)
  wire _02455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5619" *)
  wire _02456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5620" *)
  wire _02457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5620" *)
  wire _02458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5621" *)
  wire _02459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5621" *)
  wire _02460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5622" *)
  wire _02461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5622" *)
  wire _02462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5623" *)
  wire _02463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5623" *)
  wire _02464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5624" *)
  wire _02465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5624" *)
  wire _02466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5625" *)
  wire _02467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5625" *)
  wire _02468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5626" *)
  wire _02469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5626" *)
  wire _02470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5627" *)
  wire _02471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5627" *)
  wire _02472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5628" *)
  wire _02473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5628" *)
  wire _02474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5629" *)
  wire _02475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5629" *)
  wire _02476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5630" *)
  wire _02477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5630" *)
  wire _02478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5631" *)
  wire _02479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5631" *)
  wire _02480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5632" *)
  wire _02481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5632" *)
  wire _02482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5633" *)
  wire _02483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5633" *)
  wire _02484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5634" *)
  wire _02485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5634" *)
  wire _02486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5635" *)
  wire _02487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5635" *)
  wire _02488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5636" *)
  wire _02489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5636" *)
  wire _02490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5637" *)
  wire _02491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5637" *)
  wire _02492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5638" *)
  wire _02493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5638" *)
  wire _02494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5639" *)
  wire _02495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5639" *)
  wire _02496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5640" *)
  wire _02497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5640" *)
  wire _02498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5641" *)
  wire _02499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5641" *)
  wire _02500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5642" *)
  wire _02501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5642" *)
  wire _02502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5643" *)
  wire _02503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5643" *)
  wire _02504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5644" *)
  wire _02505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5644" *)
  wire _02506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5645" *)
  wire _02507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5645" *)
  wire _02508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5646" *)
  wire _02509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5646" *)
  wire _02510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5647" *)
  wire _02511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5647" *)
  wire _02512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5648" *)
  wire _02513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5648" *)
  wire _02514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5649" *)
  wire _02515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5649" *)
  wire _02516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5650" *)
  wire _02517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5650" *)
  wire _02518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5651" *)
  wire _02519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5651" *)
  wire _02520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5652" *)
  wire _02521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5652" *)
  wire _02522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5653" *)
  wire _02523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5653" *)
  wire _02524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5654" *)
  wire _02525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5654" *)
  wire _02526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5655" *)
  wire _02527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5655" *)
  wire _02528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5656" *)
  wire _02529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5656" *)
  wire _02530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5657" *)
  wire _02531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5657" *)
  wire _02532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5658" *)
  wire _02533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5658" *)
  wire _02534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5659" *)
  wire _02535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5659" *)
  wire _02536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5660" *)
  wire _02537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5660" *)
  wire _02538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5661" *)
  wire _02539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5661" *)
  wire _02540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5662" *)
  wire _02541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5662" *)
  wire _02542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5663" *)
  wire _02543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5663" *)
  wire _02544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5664" *)
  wire _02545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5664" *)
  wire _02546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5665" *)
  wire _02547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5665" *)
  wire _02548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5666" *)
  wire _02549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5666" *)
  wire _02550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5667" *)
  wire _02551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5667" *)
  wire _02552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5668" *)
  wire _02553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5668" *)
  wire _02554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5669" *)
  wire _02555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5669" *)
  wire _02556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5670" *)
  wire _02557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5670" *)
  wire _02558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5671" *)
  wire _02559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5671" *)
  wire _02560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5672" *)
  wire _02561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5672" *)
  wire _02562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5673" *)
  wire _02563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5673" *)
  wire _02564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5674" *)
  wire _02565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5674" *)
  wire _02566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5675" *)
  wire _02567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5675" *)
  wire _02568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5676" *)
  wire _02569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5676" *)
  wire _02570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5677" *)
  wire _02571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5677" *)
  wire _02572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5678" *)
  wire _02573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5678" *)
  wire _02574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5679" *)
  wire _02575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5679" *)
  wire _02576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5680" *)
  wire _02577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5680" *)
  wire _02578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5681" *)
  wire _02579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5681" *)
  wire _02580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5682" *)
  wire _02581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5682" *)
  wire _02582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5683" *)
  wire _02583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5683" *)
  wire _02584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5684" *)
  wire _02585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5684" *)
  wire _02586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5685" *)
  wire _02587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5685" *)
  wire _02588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5686" *)
  wire _02589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5686" *)
  wire _02590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5687" *)
  wire _02591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5687" *)
  wire _02592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5688" *)
  wire _02593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5688" *)
  wire _02594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5689" *)
  wire _02595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5689" *)
  wire _02596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5690" *)
  wire _02597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5690" *)
  wire _02598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5691" *)
  wire _02599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5691" *)
  wire _02600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5692" *)
  wire _02601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5692" *)
  wire _02602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5693" *)
  wire _02603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5693" *)
  wire _02604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5694" *)
  wire _02605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5694" *)
  wire _02606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5695" *)
  wire _02607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5695" *)
  wire _02608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5696" *)
  wire _02609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5696" *)
  wire _02610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5697" *)
  wire _02611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5697" *)
  wire _02612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5698" *)
  wire _02613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5698" *)
  wire _02614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5699" *)
  wire _02615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5699" *)
  wire _02616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5700" *)
  wire _02617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5700" *)
  wire _02618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5701" *)
  wire _02619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5701" *)
  wire _02620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5702" *)
  wire _02621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5702" *)
  wire _02622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5703" *)
  wire _02623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5703" *)
  wire _02624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5704" *)
  wire _02625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5704" *)
  wire _02626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5705" *)
  wire _02627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5705" *)
  wire _02628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5706" *)
  wire _02629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5706" *)
  wire _02630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5707" *)
  wire _02631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5707" *)
  wire _02632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5708" *)
  wire _02633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5708" *)
  wire _02634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5709" *)
  wire _02635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5709" *)
  wire _02636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5710" *)
  wire _02637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5710" *)
  wire _02638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5711" *)
  wire _02639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5711" *)
  wire _02640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5712" *)
  wire _02641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5712" *)
  wire _02642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5713" *)
  wire _02643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5713" *)
  wire _02644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5714" *)
  wire _02645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5714" *)
  wire _02646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5715" *)
  wire _02647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5715" *)
  wire _02648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5716" *)
  wire _02649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5716" *)
  wire _02650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5717" *)
  wire _02651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5717" *)
  wire _02652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5718" *)
  wire _02653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5718" *)
  wire _02654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5719" *)
  wire _02655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5719" *)
  wire _02656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5720" *)
  wire _02657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5720" *)
  wire _02658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5721" *)
  wire _02659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5721" *)
  wire _02660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5722" *)
  wire _02661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5722" *)
  wire _02662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5723" *)
  wire _02663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5723" *)
  wire _02664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5724" *)
  wire _02665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5724" *)
  wire _02666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5725" *)
  wire _02667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5725" *)
  wire _02668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5726" *)
  wire _02669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5726" *)
  wire _02670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5727" *)
  wire _02671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5727" *)
  wire _02672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5728" *)
  wire _02673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5728" *)
  wire _02674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5729" *)
  wire _02675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5729" *)
  wire _02676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5730" *)
  wire _02677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5730" *)
  wire _02678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5731" *)
  wire _02679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5731" *)
  wire _02680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5732" *)
  wire _02681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5732" *)
  wire _02682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5733" *)
  wire _02683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5733" *)
  wire _02684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5734" *)
  wire _02685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5734" *)
  wire _02686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5735" *)
  wire _02687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5735" *)
  wire _02688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5736" *)
  wire _02689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5736" *)
  wire _02690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5737" *)
  wire _02691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5737" *)
  wire _02692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5738" *)
  wire _02693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5738" *)
  wire _02694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5739" *)
  wire _02695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5739" *)
  wire _02696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5740" *)
  wire _02697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5740" *)
  wire _02698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5741" *)
  wire _02699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5741" *)
  wire _02700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5742" *)
  wire _02701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5742" *)
  wire _02702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5743" *)
  wire _02703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5743" *)
  wire _02704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5744" *)
  wire _02705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5744" *)
  wire _02706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5745" *)
  wire _02707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5745" *)
  wire _02708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5746" *)
  wire _02709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5746" *)
  wire _02710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5747" *)
  wire _02711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5747" *)
  wire _02712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5748" *)
  wire _02713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5748" *)
  wire _02714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5749" *)
  wire _02715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5749" *)
  wire _02716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5750" *)
  wire _02717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5750" *)
  wire _02718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5751" *)
  wire _02719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5751" *)
  wire _02720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5752" *)
  wire _02721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5752" *)
  wire _02722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5753" *)
  wire _02723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5753" *)
  wire _02724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5754" *)
  wire _02725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5754" *)
  wire _02726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5755" *)
  wire _02727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5755" *)
  wire _02728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5756" *)
  wire _02729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5756" *)
  wire _02730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5757" *)
  wire _02731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5757" *)
  wire _02732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5758" *)
  wire _02733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5758" *)
  wire _02734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5759" *)
  wire _02735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5759" *)
  wire _02736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5760" *)
  wire _02737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5760" *)
  wire _02738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5761" *)
  wire _02739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5761" *)
  wire _02740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5762" *)
  wire _02741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5762" *)
  wire _02742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5763" *)
  wire _02743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5763" *)
  wire _02744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5764" *)
  wire _02745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5764" *)
  wire _02746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5765" *)
  wire _02747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5765" *)
  wire _02748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5766" *)
  wire _02749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5766" *)
  wire _02750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5767" *)
  wire _02751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5767" *)
  wire _02752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5768" *)
  wire _02753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5768" *)
  wire _02754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5769" *)
  wire _02755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5769" *)
  wire _02756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5770" *)
  wire _02757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5770" *)
  wire _02758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5771" *)
  wire _02759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5771" *)
  wire _02760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5772" *)
  wire _02761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5772" *)
  wire _02762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5773" *)
  wire _02763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5773" *)
  wire _02764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5774" *)
  wire _02765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5774" *)
  wire _02766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5775" *)
  wire _02767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5775" *)
  wire _02768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5776" *)
  wire _02769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5776" *)
  wire _02770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5777" *)
  wire _02771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5777" *)
  wire _02772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5778" *)
  wire _02773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5778" *)
  wire _02774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5779" *)
  wire _02775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5779" *)
  wire _02776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5780" *)
  wire _02777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5780" *)
  wire _02778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5781" *)
  wire _02779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5781" *)
  wire _02780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5782" *)
  wire _02781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5782" *)
  wire _02782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5783" *)
  wire _02783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5783" *)
  wire _02784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5784" *)
  wire _02785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5784" *)
  wire _02786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5785" *)
  wire _02787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5785" *)
  wire _02788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5786" *)
  wire _02789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5786" *)
  wire _02790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5787" *)
  wire _02791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5787" *)
  wire _02792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5788" *)
  wire _02793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5788" *)
  wire _02794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5789" *)
  wire _02795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5789" *)
  wire _02796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5790" *)
  wire _02797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5790" *)
  wire _02798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5791" *)
  wire _02799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5791" *)
  wire _02800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5792" *)
  wire _02801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5792" *)
  wire _02802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5793" *)
  wire _02803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5793" *)
  wire _02804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5794" *)
  wire _02805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5794" *)
  wire _02806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5795" *)
  wire _02807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5795" *)
  wire _02808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5796" *)
  wire _02809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5796" *)
  wire _02810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5797" *)
  wire _02811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5797" *)
  wire _02812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5798" *)
  wire _02813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5798" *)
  wire _02814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5799" *)
  wire _02815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5799" *)
  wire _02816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5800" *)
  wire _02817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5800" *)
  wire _02818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5801" *)
  wire _02819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5801" *)
  wire _02820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5802" *)
  wire _02821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5802" *)
  wire _02822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5803" *)
  wire _02823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5803" *)
  wire _02824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5804" *)
  wire _02825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5804" *)
  wire _02826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5805" *)
  wire _02827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5805" *)
  wire _02828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5806" *)
  wire _02829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5806" *)
  wire _02830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5807" *)
  wire _02831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5807" *)
  wire _02832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5808" *)
  wire _02833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5808" *)
  wire _02834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5809" *)
  wire _02835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5809" *)
  wire _02836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5810" *)
  wire _02837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5810" *)
  wire _02838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5811" *)
  wire _02839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5811" *)
  wire _02840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5812" *)
  wire _02841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5812" *)
  wire _02842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5813" *)
  wire _02843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5813" *)
  wire _02844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5814" *)
  wire _02845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5814" *)
  wire _02846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5815" *)
  wire _02847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5815" *)
  wire _02848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5816" *)
  wire _02849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5816" *)
  wire _02850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5817" *)
  wire _02851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5817" *)
  wire _02852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5818" *)
  wire _02853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5818" *)
  wire _02854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5819" *)
  wire _02855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5819" *)
  wire _02856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5820" *)
  wire _02857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5820" *)
  wire _02858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5821" *)
  wire _02859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5821" *)
  wire _02860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5822" *)
  wire _02861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5822" *)
  wire _02862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5823" *)
  wire _02863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5823" *)
  wire _02864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5824" *)
  wire _02865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5824" *)
  wire _02866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5825" *)
  wire _02867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5825" *)
  wire _02868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5826" *)
  wire _02869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5826" *)
  wire _02870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5827" *)
  wire _02871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5827" *)
  wire _02872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5828" *)
  wire _02873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5828" *)
  wire _02874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5829" *)
  wire _02875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5829" *)
  wire _02876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5830" *)
  wire _02877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5830" *)
  wire _02878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5831" *)
  wire _02879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5831" *)
  wire _02880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5832" *)
  wire _02881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5832" *)
  wire _02882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5833" *)
  wire _02883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5833" *)
  wire _02884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5834" *)
  wire _02885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5834" *)
  wire _02886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5835" *)
  wire _02887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5835" *)
  wire _02888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5836" *)
  wire _02889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5836" *)
  wire _02890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5837" *)
  wire _02891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5837" *)
  wire _02892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5838" *)
  wire _02893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5838" *)
  wire _02894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5839" *)
  wire _02895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5839" *)
  wire _02896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5840" *)
  wire _02897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5840" *)
  wire _02898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5841" *)
  wire _02899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5841" *)
  wire _02900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5842" *)
  wire _02901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5842" *)
  wire _02902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5843" *)
  wire _02903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5843" *)
  wire _02904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5844" *)
  wire _02905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5844" *)
  wire _02906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5845" *)
  wire _02907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5845" *)
  wire _02908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5846" *)
  wire _02909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5846" *)
  wire _02910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5847" *)
  wire _02911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5847" *)
  wire _02912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5848" *)
  wire _02913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5848" *)
  wire _02914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5849" *)
  wire _02915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5849" *)
  wire _02916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5850" *)
  wire _02917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5850" *)
  wire _02918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5851" *)
  wire _02919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5851" *)
  wire _02920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5852" *)
  wire _02921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5852" *)
  wire _02922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5853" *)
  wire _02923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5853" *)
  wire _02924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5854" *)
  wire _02925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5854" *)
  wire _02926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5855" *)
  wire _02927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5855" *)
  wire _02928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5856" *)
  wire _02929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5856" *)
  wire _02930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5857" *)
  wire _02931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5857" *)
  wire _02932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5858" *)
  wire _02933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5858" *)
  wire _02934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5859" *)
  wire _02935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5859" *)
  wire _02936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5860" *)
  wire _02937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5860" *)
  wire _02938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5861" *)
  wire _02939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5861" *)
  wire _02940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5862" *)
  wire _02941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5862" *)
  wire _02942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5863" *)
  wire _02943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5863" *)
  wire _02944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5864" *)
  wire _02945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5864" *)
  wire _02946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5865" *)
  wire _02947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5865" *)
  wire _02948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5866" *)
  wire _02949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5866" *)
  wire _02950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5867" *)
  wire _02951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5867" *)
  wire _02952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5868" *)
  wire _02953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5868" *)
  wire _02954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5869" *)
  wire _02955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5869" *)
  wire _02956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5870" *)
  wire _02957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5870" *)
  wire _02958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5871" *)
  wire _02959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5871" *)
  wire _02960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5872" *)
  wire _02961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5872" *)
  wire _02962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5873" *)
  wire _02963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5873" *)
  wire _02964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5874" *)
  wire _02965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5874" *)
  wire _02966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5875" *)
  wire _02967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5875" *)
  wire _02968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5876" *)
  wire _02969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5876" *)
  wire _02970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5877" *)
  wire _02971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5877" *)
  wire _02972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5878" *)
  wire _02973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5878" *)
  wire _02974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5879" *)
  wire _02975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5879" *)
  wire _02976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5880" *)
  wire _02977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5880" *)
  wire _02978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5881" *)
  wire _02979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5881" *)
  wire _02980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5882" *)
  wire _02981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5882" *)
  wire _02982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5883" *)
  wire _02983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5883" *)
  wire _02984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5884" *)
  wire _02985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5884" *)
  wire _02986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5885" *)
  wire _02987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5885" *)
  wire _02988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5886" *)
  wire _02989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5886" *)
  wire _02990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5887" *)
  wire _02991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5887" *)
  wire _02992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5888" *)
  wire _02993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5888" *)
  wire _02994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5889" *)
  wire _02995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5889" *)
  wire _02996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5890" *)
  wire _02997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5890" *)
  wire _02998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5891" *)
  wire _02999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5891" *)
  wire _03000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5892" *)
  wire _03001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5892" *)
  wire _03002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5893" *)
  wire _03003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5893" *)
  wire _03004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5894" *)
  wire _03005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5894" *)
  wire _03006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5895" *)
  wire _03007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5895" *)
  wire _03008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5896" *)
  wire _03009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5896" *)
  wire _03010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5897" *)
  wire _03011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5897" *)
  wire _03012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5898" *)
  wire _03013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5898" *)
  wire _03014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5899" *)
  wire _03015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5899" *)
  wire _03016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5900" *)
  wire _03017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5900" *)
  wire _03018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5901" *)
  wire _03019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5901" *)
  wire _03020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5902" *)
  wire _03021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5902" *)
  wire _03022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5903" *)
  wire _03023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5903" *)
  wire _03024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5904" *)
  wire _03025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5904" *)
  wire _03026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5905" *)
  wire _03027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5905" *)
  wire _03028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5906" *)
  wire _03029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5906" *)
  wire _03030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5907" *)
  wire _03031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5907" *)
  wire _03032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5908" *)
  wire _03033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5908" *)
  wire _03034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5909" *)
  wire _03035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5909" *)
  wire _03036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5910" *)
  wire _03037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5910" *)
  wire _03038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5911" *)
  wire _03039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5911" *)
  wire _03040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5912" *)
  wire _03041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5912" *)
  wire _03042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5913" *)
  wire _03043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5913" *)
  wire _03044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5914" *)
  wire _03045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5914" *)
  wire _03046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5915" *)
  wire _03047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5915" *)
  wire _03048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5916" *)
  wire _03049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5916" *)
  wire _03050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5917" *)
  wire _03051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5917" *)
  wire _03052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5918" *)
  wire _03053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5918" *)
  wire _03054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5919" *)
  wire _03055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5919" *)
  wire _03056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5920" *)
  wire _03057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5920" *)
  wire _03058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5921" *)
  wire _03059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5921" *)
  wire _03060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5922" *)
  wire _03061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5922" *)
  wire _03062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5923" *)
  wire _03063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5923" *)
  wire _03064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5924" *)
  wire _03065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5924" *)
  wire _03066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5925" *)
  wire _03067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5925" *)
  wire _03068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5926" *)
  wire _03069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5926" *)
  wire _03070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5927" *)
  wire _03071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5927" *)
  wire _03072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5928" *)
  wire _03073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5928" *)
  wire _03074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5929" *)
  wire _03075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5929" *)
  wire _03076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5930" *)
  wire _03077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5930" *)
  wire _03078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5931" *)
  wire _03079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5931" *)
  wire _03080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5932" *)
  wire _03081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5932" *)
  wire _03082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5933" *)
  wire _03083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5933" *)
  wire _03084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5934" *)
  wire _03085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5934" *)
  wire _03086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5935" *)
  wire _03087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5935" *)
  wire _03088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5936" *)
  wire _03089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5936" *)
  wire _03090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5937" *)
  wire _03091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5937" *)
  wire _03092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5938" *)
  wire _03093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5938" *)
  wire _03094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5939" *)
  wire _03095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5939" *)
  wire _03096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5940" *)
  wire _03097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5940" *)
  wire _03098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5941" *)
  wire _03099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5941" *)
  wire _03100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5942" *)
  wire _03101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5942" *)
  wire _03102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5943" *)
  wire _03103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5943" *)
  wire _03104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5944" *)
  wire _03105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5944" *)
  wire _03106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5945" *)
  wire _03107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5945" *)
  wire _03108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5946" *)
  wire _03109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5946" *)
  wire _03110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5947" *)
  wire _03111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5947" *)
  wire _03112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5948" *)
  wire _03113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5948" *)
  wire _03114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5949" *)
  wire _03115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5949" *)
  wire _03116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5950" *)
  wire _03117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5950" *)
  wire _03118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5951" *)
  wire _03119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5951" *)
  wire _03120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5952" *)
  wire _03121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5952" *)
  wire _03122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5953" *)
  wire _03123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5953" *)
  wire _03124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5954" *)
  wire _03125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5954" *)
  wire _03126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5955" *)
  wire _03127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5955" *)
  wire _03128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5956" *)
  wire _03129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5956" *)
  wire _03130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5957" *)
  wire _03131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5957" *)
  wire _03132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5958" *)
  wire _03133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5958" *)
  wire _03134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5959" *)
  wire _03135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5959" *)
  wire _03136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5960" *)
  wire _03137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5960" *)
  wire _03138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5961" *)
  wire _03139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5961" *)
  wire _03140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5962" *)
  wire _03141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5962" *)
  wire _03142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5963" *)
  wire _03143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5963" *)
  wire _03144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5964" *)
  wire _03145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5964" *)
  wire _03146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5965" *)
  wire _03147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5965" *)
  wire _03148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5966" *)
  wire _03149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5966" *)
  wire _03150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5967" *)
  wire _03151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5967" *)
  wire _03152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5968" *)
  wire _03153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5968" *)
  wire _03154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5969" *)
  wire _03155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5969" *)
  wire _03156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5970" *)
  wire _03157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5970" *)
  wire _03158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5971" *)
  wire _03159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5971" *)
  wire _03160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5972" *)
  wire _03161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5972" *)
  wire _03162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5973" *)
  wire _03163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5973" *)
  wire _03164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5974" *)
  wire _03165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5974" *)
  wire _03166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5975" *)
  wire _03167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5975" *)
  wire _03168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5976" *)
  wire _03169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5976" *)
  wire _03170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5977" *)
  wire _03171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5977" *)
  wire _03172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5978" *)
  wire _03173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5978" *)
  wire _03174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5979" *)
  wire _03175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5979" *)
  wire _03176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5980" *)
  wire _03177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5980" *)
  wire _03178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5981" *)
  wire _03179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5981" *)
  wire _03180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5982" *)
  wire _03181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5982" *)
  wire _03182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5983" *)
  wire _03183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5983" *)
  wire _03184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5984" *)
  wire _03185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5984" *)
  wire _03186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5985" *)
  wire _03187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5985" *)
  wire _03188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5986" *)
  wire _03189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5986" *)
  wire _03190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5987" *)
  wire _03191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5987" *)
  wire _03192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5988" *)
  wire _03193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5988" *)
  wire _03194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5989" *)
  wire _03195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5989" *)
  wire _03196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5990" *)
  wire _03197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5990" *)
  wire _03198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5991" *)
  wire _03199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5991" *)
  wire _03200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5992" *)
  wire _03201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5992" *)
  wire _03202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5993" *)
  wire _03203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5993" *)
  wire _03204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5994" *)
  wire _03205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5994" *)
  wire _03206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5995" *)
  wire _03207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5995" *)
  wire _03208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5996" *)
  wire _03209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5996" *)
  wire _03210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5997" *)
  wire _03211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5997" *)
  wire _03212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5998" *)
  wire _03213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5998" *)
  wire _03214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5999" *)
  wire _03215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5999" *)
  wire _03216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6000" *)
  wire _03217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6000" *)
  wire _03218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6001" *)
  wire _03219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6001" *)
  wire _03220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6002" *)
  wire _03221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6002" *)
  wire _03222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6003" *)
  wire _03223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6003" *)
  wire _03224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6004" *)
  wire _03225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6004" *)
  wire _03226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6005" *)
  wire _03227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6005" *)
  wire _03228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6006" *)
  wire _03229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6006" *)
  wire _03230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6007" *)
  wire _03231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6007" *)
  wire _03232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6008" *)
  wire _03233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6008" *)
  wire _03234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6009" *)
  wire _03235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6009" *)
  wire _03236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6010" *)
  wire _03237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6010" *)
  wire _03238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6011" *)
  wire _03239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6011" *)
  wire _03240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6012" *)
  wire _03241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6012" *)
  wire _03242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6013" *)
  wire _03243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6013" *)
  wire _03244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6014" *)
  wire _03245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6014" *)
  wire _03246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6020" *)
  wire _03247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6020" *)
  wire _03248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6021" *)
  wire _03249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6021" *)
  wire _03250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6022" *)
  wire _03251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6022" *)
  wire _03252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6023" *)
  wire _03253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6023" *)
  wire _03254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6024" *)
  wire _03255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6024" *)
  wire _03256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6025" *)
  wire _03257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6025" *)
  wire _03258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6026" *)
  wire _03259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6026" *)
  wire _03260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6027" *)
  wire _03261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6027" *)
  wire _03262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6028" *)
  wire _03263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6028" *)
  wire _03264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6029" *)
  wire _03265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6029" *)
  wire _03266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6030" *)
  wire _03267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6030" *)
  wire _03268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6031" *)
  wire _03269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6031" *)
  wire _03270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6032" *)
  wire _03271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6032" *)
  wire _03272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6033" *)
  wire _03273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6033" *)
  wire _03274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6034" *)
  wire _03275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6034" *)
  wire _03276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6035" *)
  wire _03277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6035" *)
  wire _03278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6036" *)
  wire _03279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6036" *)
  wire _03280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6037" *)
  wire _03281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6037" *)
  wire _03282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6038" *)
  wire _03283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6038" *)
  wire _03284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6039" *)
  wire _03285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6039" *)
  wire _03286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6040" *)
  wire _03287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6040" *)
  wire _03288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6041" *)
  wire _03289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6041" *)
  wire _03290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6042" *)
  wire _03291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6042" *)
  wire _03292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6043" *)
  wire _03293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6043" *)
  wire _03294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6044" *)
  wire _03295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6044" *)
  wire _03296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6045" *)
  wire _03297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6045" *)
  wire _03298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6046" *)
  wire _03299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6046" *)
  wire _03300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6047" *)
  wire _03301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6047" *)
  wire _03302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6048" *)
  wire _03303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6048" *)
  wire _03304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6049" *)
  wire _03305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6049" *)
  wire _03306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6050" *)
  wire _03307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6050" *)
  wire _03308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6051" *)
  wire _03309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6051" *)
  wire _03310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6052" *)
  wire _03311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6052" *)
  wire _03312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6053" *)
  wire _03313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6053" *)
  wire _03314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6054" *)
  wire _03315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6054" *)
  wire _03316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6055" *)
  wire _03317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6055" *)
  wire _03318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6056" *)
  wire _03319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6056" *)
  wire _03320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6057" *)
  wire _03321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6057" *)
  wire _03322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6058" *)
  wire _03323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6058" *)
  wire _03324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6059" *)
  wire _03325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6059" *)
  wire _03326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6060" *)
  wire _03327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6060" *)
  wire _03328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6061" *)
  wire _03329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6061" *)
  wire _03330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6062" *)
  wire _03331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6062" *)
  wire _03332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6063" *)
  wire _03333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6063" *)
  wire _03334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6064" *)
  wire _03335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6064" *)
  wire _03336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6065" *)
  wire _03337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6065" *)
  wire _03338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6066" *)
  wire _03339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6066" *)
  wire _03340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6067" *)
  wire _03341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6067" *)
  wire _03342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6068" *)
  wire _03343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6068" *)
  wire _03344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6069" *)
  wire _03345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6069" *)
  wire _03346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6070" *)
  wire _03347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6070" *)
  wire _03348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6071" *)
  wire _03349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6071" *)
  wire _03350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6072" *)
  wire _03351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6072" *)
  wire _03352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6073" *)
  wire _03353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6073" *)
  wire _03354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6074" *)
  wire _03355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6074" *)
  wire _03356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6075" *)
  wire _03357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6075" *)
  wire _03358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6076" *)
  wire _03359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6076" *)
  wire _03360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6077" *)
  wire _03361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6077" *)
  wire _03362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6078" *)
  wire _03363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6078" *)
  wire _03364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6079" *)
  wire _03365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6079" *)
  wire _03366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6080" *)
  wire _03367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6080" *)
  wire _03368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6081" *)
  wire _03369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6081" *)
  wire _03370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6082" *)
  wire _03371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6082" *)
  wire _03372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6083" *)
  wire _03373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6083" *)
  wire _03374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6084" *)
  wire _03375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6084" *)
  wire _03376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6085" *)
  wire _03377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6085" *)
  wire _03378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6086" *)
  wire _03379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6086" *)
  wire _03380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6087" *)
  wire _03381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6087" *)
  wire _03382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6088" *)
  wire _03383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6088" *)
  wire _03384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6089" *)
  wire _03385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6089" *)
  wire _03386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6090" *)
  wire _03387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6090" *)
  wire _03388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6091" *)
  wire _03389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6091" *)
  wire _03390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6092" *)
  wire _03391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6092" *)
  wire _03392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6093" *)
  wire _03393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6093" *)
  wire _03394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6094" *)
  wire _03395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6094" *)
  wire _03396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6095" *)
  wire _03397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6095" *)
  wire _03398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6096" *)
  wire _03399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6096" *)
  wire _03400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6097" *)
  wire _03401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6097" *)
  wire _03402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6098" *)
  wire _03403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6098" *)
  wire _03404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6099" *)
  wire _03405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6099" *)
  wire _03406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6100" *)
  wire _03407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6100" *)
  wire _03408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6101" *)
  wire _03409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6101" *)
  wire _03410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6102" *)
  wire _03411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6102" *)
  wire _03412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6103" *)
  wire _03413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6103" *)
  wire _03414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6104" *)
  wire _03415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6104" *)
  wire _03416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6105" *)
  wire _03417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6105" *)
  wire _03418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6106" *)
  wire _03419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6106" *)
  wire _03420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6107" *)
  wire _03421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6107" *)
  wire _03422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6108" *)
  wire _03423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6108" *)
  wire _03424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6109" *)
  wire _03425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6109" *)
  wire _03426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6110" *)
  wire _03427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6110" *)
  wire _03428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6111" *)
  wire _03429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6111" *)
  wire _03430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6112" *)
  wire _03431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6112" *)
  wire _03432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6113" *)
  wire _03433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6113" *)
  wire _03434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6114" *)
  wire _03435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6114" *)
  wire _03436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6115" *)
  wire _03437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6115" *)
  wire _03438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6116" *)
  wire _03439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6116" *)
  wire _03440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6117" *)
  wire _03441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6117" *)
  wire _03442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6118" *)
  wire _03443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6118" *)
  wire _03444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6119" *)
  wire _03445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6119" *)
  wire _03446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6120" *)
  wire _03447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6120" *)
  wire _03448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6121" *)
  wire _03449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6121" *)
  wire _03450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6122" *)
  wire _03451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6122" *)
  wire _03452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6123" *)
  wire _03453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6123" *)
  wire _03454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6124" *)
  wire _03455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6124" *)
  wire _03456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6125" *)
  wire _03457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6125" *)
  wire _03458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6126" *)
  wire _03459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6126" *)
  wire _03460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6127" *)
  wire _03461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6127" *)
  wire _03462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6128" *)
  wire _03463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6128" *)
  wire _03464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6129" *)
  wire _03465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6129" *)
  wire _03466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6130" *)
  wire _03467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6130" *)
  wire _03468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6131" *)
  wire _03469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6131" *)
  wire _03470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6132" *)
  wire _03471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6132" *)
  wire _03472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6133" *)
  wire _03473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6133" *)
  wire _03474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6134" *)
  wire _03475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6134" *)
  wire _03476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6135" *)
  wire _03477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6135" *)
  wire _03478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6136" *)
  wire _03479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6136" *)
  wire _03480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6137" *)
  wire _03481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6137" *)
  wire _03482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6138" *)
  wire _03483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6138" *)
  wire _03484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6139" *)
  wire _03485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6139" *)
  wire _03486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6140" *)
  wire _03487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6140" *)
  wire _03488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6141" *)
  wire _03489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6141" *)
  wire _03490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6142" *)
  wire _03491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6142" *)
  wire _03492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6143" *)
  wire _03493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6143" *)
  wire _03494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6144" *)
  wire _03495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6144" *)
  wire _03496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6145" *)
  wire _03497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6145" *)
  wire _03498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6146" *)
  wire _03499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6146" *)
  wire _03500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6147" *)
  wire _03501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6147" *)
  wire _03502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6148" *)
  wire _03503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6148" *)
  wire _03504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6149" *)
  wire _03505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6149" *)
  wire _03506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6150" *)
  wire _03507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6150" *)
  wire _03508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6151" *)
  wire _03509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6151" *)
  wire _03510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6152" *)
  wire _03511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6152" *)
  wire _03512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6153" *)
  wire _03513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6153" *)
  wire _03514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6154" *)
  wire _03515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6154" *)
  wire _03516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6155" *)
  wire _03517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6155" *)
  wire _03518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6156" *)
  wire _03519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6156" *)
  wire _03520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6157" *)
  wire _03521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6157" *)
  wire _03522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6158" *)
  wire _03523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6158" *)
  wire _03524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6159" *)
  wire _03525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6159" *)
  wire _03526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6160" *)
  wire _03527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6160" *)
  wire _03528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6161" *)
  wire _03529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6161" *)
  wire _03530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6162" *)
  wire _03531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6162" *)
  wire _03532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6163" *)
  wire _03533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6163" *)
  wire _03534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6164" *)
  wire _03535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6164" *)
  wire _03536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6165" *)
  wire _03537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6165" *)
  wire _03538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6166" *)
  wire _03539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6166" *)
  wire _03540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6167" *)
  wire _03541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6167" *)
  wire _03542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6168" *)
  wire _03543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6168" *)
  wire _03544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6169" *)
  wire _03545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6169" *)
  wire _03546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6170" *)
  wire _03547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6170" *)
  wire _03548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6171" *)
  wire _03549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6171" *)
  wire _03550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6172" *)
  wire _03551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6172" *)
  wire _03552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6173" *)
  wire _03553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6173" *)
  wire _03554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6174" *)
  wire _03555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6174" *)
  wire _03556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6175" *)
  wire _03557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6175" *)
  wire _03558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6176" *)
  wire _03559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6176" *)
  wire _03560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6177" *)
  wire _03561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6177" *)
  wire _03562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6178" *)
  wire _03563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6178" *)
  wire _03564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6179" *)
  wire _03565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6179" *)
  wire _03566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6180" *)
  wire _03567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6180" *)
  wire _03568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6181" *)
  wire _03569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6181" *)
  wire _03570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6182" *)
  wire _03571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6182" *)
  wire _03572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6183" *)
  wire _03573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6183" *)
  wire _03574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6184" *)
  wire _03575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6184" *)
  wire _03576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6185" *)
  wire _03577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6185" *)
  wire _03578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6186" *)
  wire _03579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6186" *)
  wire _03580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6187" *)
  wire _03581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6187" *)
  wire _03582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6188" *)
  wire _03583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6188" *)
  wire _03584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6189" *)
  wire _03585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6189" *)
  wire _03586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6190" *)
  wire _03587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6190" *)
  wire _03588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6191" *)
  wire _03589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6191" *)
  wire _03590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6192" *)
  wire _03591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6192" *)
  wire _03592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6193" *)
  wire _03593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6193" *)
  wire _03594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6194" *)
  wire _03595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6194" *)
  wire _03596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6195" *)
  wire _03597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6195" *)
  wire _03598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6196" *)
  wire _03599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6196" *)
  wire _03600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6197" *)
  wire _03601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6197" *)
  wire _03602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6198" *)
  wire _03603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6198" *)
  wire _03604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6199" *)
  wire _03605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6199" *)
  wire _03606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6200" *)
  wire _03607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6200" *)
  wire _03608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6201" *)
  wire _03609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6201" *)
  wire _03610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6202" *)
  wire _03611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6202" *)
  wire _03612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6203" *)
  wire _03613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6203" *)
  wire _03614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6204" *)
  wire _03615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6204" *)
  wire _03616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6205" *)
  wire _03617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6205" *)
  wire _03618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6206" *)
  wire _03619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6206" *)
  wire _03620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6207" *)
  wire _03621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6207" *)
  wire _03622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6208" *)
  wire _03623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6208" *)
  wire _03624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6209" *)
  wire _03625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6209" *)
  wire _03626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6210" *)
  wire _03627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6210" *)
  wire _03628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6211" *)
  wire _03629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6211" *)
  wire _03630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6212" *)
  wire _03631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6212" *)
  wire _03632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6213" *)
  wire _03633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6213" *)
  wire _03634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6214" *)
  wire _03635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6214" *)
  wire _03636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6215" *)
  wire _03637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6215" *)
  wire _03638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6216" *)
  wire _03639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6216" *)
  wire _03640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6217" *)
  wire _03641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6217" *)
  wire _03642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6218" *)
  wire _03643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6218" *)
  wire _03644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6219" *)
  wire _03645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6219" *)
  wire _03646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6220" *)
  wire _03647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6220" *)
  wire _03648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6221" *)
  wire _03649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6221" *)
  wire _03650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6222" *)
  wire _03651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6222" *)
  wire _03652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6223" *)
  wire _03653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6223" *)
  wire _03654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6224" *)
  wire _03655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6224" *)
  wire _03656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6225" *)
  wire _03657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6225" *)
  wire _03658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6226" *)
  wire _03659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6226" *)
  wire _03660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6227" *)
  wire _03661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6227" *)
  wire _03662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6228" *)
  wire _03663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6228" *)
  wire _03664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6229" *)
  wire _03665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6229" *)
  wire _03666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6230" *)
  wire _03667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6230" *)
  wire _03668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6231" *)
  wire _03669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6231" *)
  wire _03670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6232" *)
  wire _03671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6232" *)
  wire _03672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6233" *)
  wire _03673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6233" *)
  wire _03674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6234" *)
  wire _03675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6234" *)
  wire _03676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6235" *)
  wire _03677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6235" *)
  wire _03678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6236" *)
  wire _03679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6236" *)
  wire _03680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6237" *)
  wire _03681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6237" *)
  wire _03682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6238" *)
  wire _03683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6238" *)
  wire _03684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6239" *)
  wire _03685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6239" *)
  wire _03686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6240" *)
  wire _03687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6240" *)
  wire _03688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6241" *)
  wire _03689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6241" *)
  wire _03690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6242" *)
  wire _03691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6242" *)
  wire _03692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6243" *)
  wire _03693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6243" *)
  wire _03694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6244" *)
  wire _03695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6244" *)
  wire _03696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6245" *)
  wire _03697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6245" *)
  wire _03698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6246" *)
  wire _03699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6246" *)
  wire _03700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6247" *)
  wire _03701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6247" *)
  wire _03702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6248" *)
  wire _03703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6248" *)
  wire _03704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6249" *)
  wire _03705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6249" *)
  wire _03706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6250" *)
  wire _03707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6250" *)
  wire _03708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6251" *)
  wire _03709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6251" *)
  wire _03710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6252" *)
  wire _03711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6252" *)
  wire _03712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6253" *)
  wire _03713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6253" *)
  wire _03714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6254" *)
  wire _03715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6254" *)
  wire _03716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6255" *)
  wire _03717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6255" *)
  wire _03718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6256" *)
  wire _03719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6256" *)
  wire _03720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6257" *)
  wire _03721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6257" *)
  wire _03722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6258" *)
  wire _03723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6258" *)
  wire _03724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6259" *)
  wire _03725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6259" *)
  wire _03726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6260" *)
  wire _03727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6260" *)
  wire _03728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6261" *)
  wire _03729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6261" *)
  wire _03730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6262" *)
  wire _03731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6262" *)
  wire _03732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6263" *)
  wire _03733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6263" *)
  wire _03734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6264" *)
  wire _03735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6264" *)
  wire _03736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6265" *)
  wire _03737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6265" *)
  wire _03738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6266" *)
  wire _03739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6266" *)
  wire _03740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6267" *)
  wire _03741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6267" *)
  wire _03742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6268" *)
  wire _03743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6268" *)
  wire _03744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6269" *)
  wire _03745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6269" *)
  wire _03746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6270" *)
  wire _03747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6270" *)
  wire _03748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6271" *)
  wire _03749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6271" *)
  wire _03750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6272" *)
  wire _03751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6272" *)
  wire _03752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6273" *)
  wire _03753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6273" *)
  wire _03754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6274" *)
  wire _03755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6274" *)
  wire _03756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6275" *)
  wire _03757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6275" *)
  wire _03758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6276" *)
  wire _03759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6276" *)
  wire _03760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6277" *)
  wire _03761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6277" *)
  wire _03762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6278" *)
  wire _03763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6278" *)
  wire _03764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6279" *)
  wire _03765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6279" *)
  wire _03766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6280" *)
  wire _03767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6280" *)
  wire _03768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6281" *)
  wire _03769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6281" *)
  wire _03770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6282" *)
  wire _03771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6282" *)
  wire _03772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6283" *)
  wire _03773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6283" *)
  wire _03774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6284" *)
  wire _03775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6284" *)
  wire _03776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6285" *)
  wire _03777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6285" *)
  wire _03778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6286" *)
  wire _03779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6286" *)
  wire _03780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6287" *)
  wire _03781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6287" *)
  wire _03782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6288" *)
  wire _03783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6288" *)
  wire _03784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6289" *)
  wire _03785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6289" *)
  wire _03786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6290" *)
  wire _03787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6290" *)
  wire _03788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6291" *)
  wire _03789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6291" *)
  wire _03790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6292" *)
  wire _03791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6292" *)
  wire _03792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6293" *)
  wire _03793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6293" *)
  wire _03794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6294" *)
  wire _03795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6294" *)
  wire _03796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6295" *)
  wire _03797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6295" *)
  wire _03798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6296" *)
  wire _03799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6296" *)
  wire _03800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6297" *)
  wire _03801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6297" *)
  wire _03802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6298" *)
  wire _03803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6298" *)
  wire _03804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6299" *)
  wire _03805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6299" *)
  wire _03806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6300" *)
  wire _03807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6300" *)
  wire _03808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6301" *)
  wire _03809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6301" *)
  wire _03810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6302" *)
  wire _03811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6302" *)
  wire _03812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6303" *)
  wire _03813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6303" *)
  wire _03814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6304" *)
  wire _03815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6304" *)
  wire _03816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6305" *)
  wire _03817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6305" *)
  wire _03818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6306" *)
  wire _03819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6306" *)
  wire _03820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6307" *)
  wire _03821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6307" *)
  wire _03822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6308" *)
  wire _03823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6308" *)
  wire _03824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6309" *)
  wire _03825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6309" *)
  wire _03826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6310" *)
  wire _03827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6310" *)
  wire _03828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6311" *)
  wire _03829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6311" *)
  wire _03830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6312" *)
  wire _03831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6312" *)
  wire _03832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6313" *)
  wire _03833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6313" *)
  wire _03834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6314" *)
  wire _03835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6314" *)
  wire _03836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6315" *)
  wire _03837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6315" *)
  wire _03838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6316" *)
  wire _03839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6316" *)
  wire _03840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6317" *)
  wire _03841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6317" *)
  wire _03842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6318" *)
  wire _03843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6318" *)
  wire _03844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6319" *)
  wire _03845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6319" *)
  wire _03846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6320" *)
  wire _03847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6320" *)
  wire _03848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6321" *)
  wire _03849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6321" *)
  wire _03850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6322" *)
  wire _03851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6322" *)
  wire _03852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6323" *)
  wire _03853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6323" *)
  wire _03854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6324" *)
  wire _03855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6324" *)
  wire _03856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6325" *)
  wire _03857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6325" *)
  wire _03858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6326" *)
  wire _03859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6326" *)
  wire _03860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6327" *)
  wire _03861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6327" *)
  wire _03862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6328" *)
  wire _03863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6328" *)
  wire _03864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6329" *)
  wire _03865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6329" *)
  wire _03866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6330" *)
  wire _03867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6330" *)
  wire _03868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6331" *)
  wire _03869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6331" *)
  wire _03870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6332" *)
  wire _03871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6332" *)
  wire _03872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6333" *)
  wire _03873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6333" *)
  wire _03874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6334" *)
  wire _03875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6334" *)
  wire _03876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6335" *)
  wire _03877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6335" *)
  wire _03878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6336" *)
  wire _03879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6336" *)
  wire _03880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6337" *)
  wire _03881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6337" *)
  wire _03882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6338" *)
  wire _03883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6338" *)
  wire _03884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6339" *)
  wire _03885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6339" *)
  wire _03886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6340" *)
  wire _03887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6340" *)
  wire _03888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6341" *)
  wire _03889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6341" *)
  wire _03890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6342" *)
  wire _03891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6342" *)
  wire _03892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6343" *)
  wire _03893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6343" *)
  wire _03894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6344" *)
  wire _03895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6344" *)
  wire _03896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6345" *)
  wire _03897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6345" *)
  wire _03898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6346" *)
  wire _03899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6346" *)
  wire _03900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6347" *)
  wire _03901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6347" *)
  wire _03902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6348" *)
  wire _03903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6348" *)
  wire _03904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6349" *)
  wire _03905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6349" *)
  wire _03906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6350" *)
  wire _03907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6350" *)
  wire _03908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6351" *)
  wire _03909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6351" *)
  wire _03910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6352" *)
  wire _03911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6352" *)
  wire _03912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6353" *)
  wire _03913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6353" *)
  wire _03914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6354" *)
  wire _03915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6354" *)
  wire _03916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6355" *)
  wire _03917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6355" *)
  wire _03918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6356" *)
  wire _03919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6356" *)
  wire _03920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6357" *)
  wire _03921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6357" *)
  wire _03922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6358" *)
  wire _03923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6358" *)
  wire _03924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6359" *)
  wire _03925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6359" *)
  wire _03926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6360" *)
  wire _03927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6360" *)
  wire _03928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6361" *)
  wire _03929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6361" *)
  wire _03930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6362" *)
  wire _03931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6362" *)
  wire _03932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6363" *)
  wire _03933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6363" *)
  wire _03934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6364" *)
  wire _03935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6364" *)
  wire _03936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6365" *)
  wire _03937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6365" *)
  wire _03938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6366" *)
  wire _03939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6366" *)
  wire _03940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6367" *)
  wire _03941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6367" *)
  wire _03942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6368" *)
  wire _03943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6368" *)
  wire _03944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6369" *)
  wire _03945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6369" *)
  wire _03946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6370" *)
  wire _03947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6370" *)
  wire _03948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6371" *)
  wire _03949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6371" *)
  wire _03950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6372" *)
  wire _03951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6372" *)
  wire _03952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6373" *)
  wire _03953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6373" *)
  wire _03954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6374" *)
  wire _03955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6374" *)
  wire _03956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6375" *)
  wire _03957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6375" *)
  wire _03958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6376" *)
  wire _03959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6376" *)
  wire _03960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6377" *)
  wire _03961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6377" *)
  wire _03962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6378" *)
  wire _03963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6378" *)
  wire _03964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6379" *)
  wire _03965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6379" *)
  wire _03966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6380" *)
  wire _03967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6380" *)
  wire _03968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6381" *)
  wire _03969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6381" *)
  wire _03970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6382" *)
  wire _03971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6382" *)
  wire _03972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6383" *)
  wire _03973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6383" *)
  wire _03974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6384" *)
  wire _03975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6384" *)
  wire _03976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6385" *)
  wire _03977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6385" *)
  wire _03978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6386" *)
  wire _03979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6386" *)
  wire _03980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6387" *)
  wire _03981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6387" *)
  wire _03982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6388" *)
  wire _03983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6388" *)
  wire _03984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6389" *)
  wire _03985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6389" *)
  wire _03986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6390" *)
  wire _03987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6390" *)
  wire _03988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6391" *)
  wire _03989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6391" *)
  wire _03990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6392" *)
  wire _03991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6392" *)
  wire _03992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6393" *)
  wire _03993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6393" *)
  wire _03994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6394" *)
  wire _03995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6394" *)
  wire _03996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6395" *)
  wire _03997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6395" *)
  wire _03998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6396" *)
  wire _03999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6396" *)
  wire _04000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6397" *)
  wire _04001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6397" *)
  wire _04002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6398" *)
  wire _04003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6398" *)
  wire _04004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6399" *)
  wire _04005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6399" *)
  wire _04006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6400" *)
  wire _04007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6400" *)
  wire _04008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6401" *)
  wire _04009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6401" *)
  wire _04010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6402" *)
  wire _04011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6402" *)
  wire _04012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6403" *)
  wire _04013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6403" *)
  wire _04014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6404" *)
  wire _04015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6404" *)
  wire _04016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6405" *)
  wire _04017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6405" *)
  wire _04018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6406" *)
  wire _04019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6406" *)
  wire _04020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6407" *)
  wire _04021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6407" *)
  wire _04022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6408" *)
  wire _04023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6408" *)
  wire _04024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6409" *)
  wire _04025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6409" *)
  wire _04026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6410" *)
  wire _04027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6410" *)
  wire _04028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6411" *)
  wire _04029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6411" *)
  wire _04030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6412" *)
  wire _04031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6412" *)
  wire _04032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6413" *)
  wire _04033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6413" *)
  wire _04034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6414" *)
  wire _04035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6414" *)
  wire _04036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6415" *)
  wire _04037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6415" *)
  wire _04038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6416" *)
  wire _04039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6416" *)
  wire _04040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6417" *)
  wire _04041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6417" *)
  wire _04042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6418" *)
  wire _04043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6418" *)
  wire _04044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6419" *)
  wire _04045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6419" *)
  wire _04046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6420" *)
  wire _04047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6420" *)
  wire _04048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6421" *)
  wire _04049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6421" *)
  wire _04050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6422" *)
  wire _04051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6422" *)
  wire _04052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6423" *)
  wire _04053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6423" *)
  wire _04054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6424" *)
  wire _04055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6424" *)
  wire _04056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6425" *)
  wire _04057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6425" *)
  wire _04058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6426" *)
  wire _04059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6426" *)
  wire _04060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6427" *)
  wire _04061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6427" *)
  wire _04062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6428" *)
  wire _04063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6428" *)
  wire _04064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6429" *)
  wire _04065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6429" *)
  wire _04066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6430" *)
  wire _04067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6430" *)
  wire _04068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6431" *)
  wire _04069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6431" *)
  wire _04070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6432" *)
  wire _04071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6432" *)
  wire _04072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6433" *)
  wire _04073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6433" *)
  wire _04074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6434" *)
  wire _04075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6434" *)
  wire _04076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6435" *)
  wire _04077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6435" *)
  wire _04078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6436" *)
  wire _04079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6436" *)
  wire _04080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6437" *)
  wire _04081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6437" *)
  wire _04082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6438" *)
  wire _04083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6438" *)
  wire _04084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6439" *)
  wire _04085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6439" *)
  wire _04086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6440" *)
  wire _04087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6440" *)
  wire _04088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6441" *)
  wire _04089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6441" *)
  wire _04090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6442" *)
  wire _04091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6442" *)
  wire _04092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6443" *)
  wire _04093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6443" *)
  wire _04094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6444" *)
  wire _04095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6444" *)
  wire _04096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6445" *)
  wire _04097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6445" *)
  wire _04098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6446" *)
  wire _04099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6446" *)
  wire _04100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6447" *)
  wire _04101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6447" *)
  wire _04102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6448" *)
  wire _04103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6448" *)
  wire _04104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6449" *)
  wire _04105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6449" *)
  wire _04106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6450" *)
  wire _04107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6450" *)
  wire _04108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6451" *)
  wire _04109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6451" *)
  wire _04110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6452" *)
  wire _04111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6452" *)
  wire _04112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6453" *)
  wire _04113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6453" *)
  wire _04114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6454" *)
  wire _04115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6454" *)
  wire _04116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6455" *)
  wire _04117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6455" *)
  wire _04118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6456" *)
  wire _04119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6456" *)
  wire _04120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6457" *)
  wire _04121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6457" *)
  wire _04122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6458" *)
  wire _04123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6458" *)
  wire _04124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6459" *)
  wire _04125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6459" *)
  wire _04126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6460" *)
  wire _04127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6460" *)
  wire _04128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6461" *)
  wire _04129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6461" *)
  wire _04130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6462" *)
  wire _04131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6462" *)
  wire _04132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6463" *)
  wire _04133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6463" *)
  wire _04134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6464" *)
  wire _04135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6464" *)
  wire _04136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6465" *)
  wire _04137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6465" *)
  wire _04138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6466" *)
  wire _04139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6466" *)
  wire _04140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6467" *)
  wire _04141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6467" *)
  wire _04142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6468" *)
  wire _04143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6468" *)
  wire _04144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6469" *)
  wire _04145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6469" *)
  wire _04146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6470" *)
  wire _04147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6470" *)
  wire _04148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6471" *)
  wire _04149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6471" *)
  wire _04150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6472" *)
  wire _04151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6472" *)
  wire _04152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6473" *)
  wire _04153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6473" *)
  wire _04154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6474" *)
  wire _04155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6474" *)
  wire _04156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6475" *)
  wire _04157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6475" *)
  wire _04158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6476" *)
  wire _04159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6476" *)
  wire _04160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6477" *)
  wire _04161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6477" *)
  wire _04162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6478" *)
  wire _04163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6478" *)
  wire _04164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6479" *)
  wire _04165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6479" *)
  wire _04166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6480" *)
  wire _04167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6480" *)
  wire _04168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6481" *)
  wire _04169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6481" *)
  wire _04170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6482" *)
  wire _04171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6482" *)
  wire _04172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6483" *)
  wire _04173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6483" *)
  wire _04174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6484" *)
  wire _04175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6484" *)
  wire _04176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6485" *)
  wire _04177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6485" *)
  wire _04178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6486" *)
  wire _04179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6486" *)
  wire _04180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6487" *)
  wire _04181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6487" *)
  wire _04182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6488" *)
  wire _04183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6488" *)
  wire _04184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6489" *)
  wire _04185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6489" *)
  wire _04186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6490" *)
  wire _04187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6490" *)
  wire _04188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6491" *)
  wire _04189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6491" *)
  wire _04190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6492" *)
  wire _04191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6492" *)
  wire _04192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6493" *)
  wire _04193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6493" *)
  wire _04194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6494" *)
  wire _04195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6494" *)
  wire _04196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6495" *)
  wire _04197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6495" *)
  wire _04198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6496" *)
  wire _04199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6496" *)
  wire _04200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6497" *)
  wire _04201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6497" *)
  wire _04202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6498" *)
  wire _04203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6498" *)
  wire _04204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6499" *)
  wire _04205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6499" *)
  wire _04206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6500" *)
  wire _04207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6500" *)
  wire _04208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6501" *)
  wire _04209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6501" *)
  wire _04210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6502" *)
  wire _04211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6502" *)
  wire _04212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6503" *)
  wire _04213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6503" *)
  wire _04214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6504" *)
  wire _04215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6504" *)
  wire _04216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6505" *)
  wire _04217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6505" *)
  wire _04218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6506" *)
  wire _04219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6506" *)
  wire _04220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6507" *)
  wire _04221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6507" *)
  wire _04222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6508" *)
  wire _04223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6508" *)
  wire _04224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6509" *)
  wire _04225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6509" *)
  wire _04226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6510" *)
  wire _04227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6510" *)
  wire _04228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6511" *)
  wire _04229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6511" *)
  wire _04230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6512" *)
  wire _04231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6512" *)
  wire _04232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6513" *)
  wire _04233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6513" *)
  wire _04234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6514" *)
  wire _04235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6514" *)
  wire _04236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6515" *)
  wire _04237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6515" *)
  wire _04238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6516" *)
  wire _04239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6516" *)
  wire _04240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6517" *)
  wire _04241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6517" *)
  wire _04242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6518" *)
  wire _04243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6518" *)
  wire _04244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6519" *)
  wire _04245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6519" *)
  wire _04246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6520" *)
  wire _04247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6520" *)
  wire _04248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6521" *)
  wire _04249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6521" *)
  wire _04250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6522" *)
  wire _04251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6522" *)
  wire _04252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6523" *)
  wire _04253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6523" *)
  wire _04254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6524" *)
  wire _04255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6524" *)
  wire _04256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6525" *)
  wire _04257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6525" *)
  wire _04258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6526" *)
  wire _04259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6526" *)
  wire _04260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6527" *)
  wire _04261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6527" *)
  wire _04262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6528" *)
  wire _04263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6528" *)
  wire _04264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6529" *)
  wire _04265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6529" *)
  wire _04266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6530" *)
  wire _04267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6530" *)
  wire _04268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6536" *)
  wire _04269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6536" *)
  wire _04270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6537" *)
  wire _04271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6537" *)
  wire _04272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6538" *)
  wire _04273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6538" *)
  wire _04274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6539" *)
  wire _04275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6539" *)
  wire _04276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6540" *)
  wire _04277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6540" *)
  wire _04278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6541" *)
  wire _04279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6541" *)
  wire _04280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6542" *)
  wire _04281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6542" *)
  wire _04282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6543" *)
  wire _04283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6543" *)
  wire _04284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6544" *)
  wire _04285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6544" *)
  wire _04286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6545" *)
  wire _04287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6545" *)
  wire _04288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6546" *)
  wire _04289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6546" *)
  wire _04290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6547" *)
  wire _04291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6547" *)
  wire _04292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6548" *)
  wire _04293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6548" *)
  wire _04294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6549" *)
  wire _04295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6549" *)
  wire _04296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6550" *)
  wire _04297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6550" *)
  wire _04298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6551" *)
  wire _04299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6551" *)
  wire _04300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6552" *)
  wire _04301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6552" *)
  wire _04302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6553" *)
  wire _04303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6553" *)
  wire _04304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6554" *)
  wire _04305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6554" *)
  wire _04306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6555" *)
  wire _04307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6555" *)
  wire _04308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6556" *)
  wire _04309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6556" *)
  wire _04310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6557" *)
  wire _04311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6557" *)
  wire _04312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6558" *)
  wire _04313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6558" *)
  wire _04314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6559" *)
  wire _04315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6559" *)
  wire _04316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6560" *)
  wire _04317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6560" *)
  wire _04318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6561" *)
  wire _04319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6561" *)
  wire _04320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6562" *)
  wire _04321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6562" *)
  wire _04322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6563" *)
  wire _04323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6563" *)
  wire _04324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6564" *)
  wire _04325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6564" *)
  wire _04326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6565" *)
  wire _04327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6565" *)
  wire _04328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6566" *)
  wire _04329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6566" *)
  wire _04330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6567" *)
  wire _04331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6567" *)
  wire _04332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6568" *)
  wire _04333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6568" *)
  wire _04334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6569" *)
  wire _04335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6569" *)
  wire _04336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6570" *)
  wire _04337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6570" *)
  wire _04338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6571" *)
  wire _04339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6571" *)
  wire _04340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6572" *)
  wire _04341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6572" *)
  wire _04342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6573" *)
  wire _04343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6573" *)
  wire _04344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6574" *)
  wire _04345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6574" *)
  wire _04346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6575" *)
  wire _04347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6575" *)
  wire _04348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6576" *)
  wire _04349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6576" *)
  wire _04350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6577" *)
  wire _04351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6577" *)
  wire _04352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6578" *)
  wire _04353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6578" *)
  wire _04354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6579" *)
  wire _04355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6579" *)
  wire _04356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6580" *)
  wire _04357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6580" *)
  wire _04358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6581" *)
  wire _04359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6581" *)
  wire _04360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6582" *)
  wire _04361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6582" *)
  wire _04362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6583" *)
  wire _04363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6583" *)
  wire _04364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6584" *)
  wire _04365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6584" *)
  wire _04366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6585" *)
  wire _04367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6585" *)
  wire _04368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6586" *)
  wire _04369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6586" *)
  wire _04370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6587" *)
  wire _04371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6587" *)
  wire _04372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6588" *)
  wire _04373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6588" *)
  wire _04374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6589" *)
  wire _04375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6589" *)
  wire _04376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6590" *)
  wire _04377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6590" *)
  wire _04378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6591" *)
  wire _04379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6591" *)
  wire _04380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6592" *)
  wire _04381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6592" *)
  wire _04382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6593" *)
  wire _04383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6593" *)
  wire _04384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6594" *)
  wire _04385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6594" *)
  wire _04386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6595" *)
  wire _04387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6595" *)
  wire _04388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6596" *)
  wire _04389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6596" *)
  wire _04390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6597" *)
  wire _04391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6597" *)
  wire _04392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6598" *)
  wire _04393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6598" *)
  wire _04394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6599" *)
  wire _04395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6599" *)
  wire _04396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6600" *)
  wire _04397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6600" *)
  wire _04398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6601" *)
  wire _04399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6601" *)
  wire _04400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6602" *)
  wire _04401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6602" *)
  wire _04402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6603" *)
  wire _04403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6603" *)
  wire _04404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6604" *)
  wire _04405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6604" *)
  wire _04406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6605" *)
  wire _04407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6605" *)
  wire _04408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6606" *)
  wire _04409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6606" *)
  wire _04410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6607" *)
  wire _04411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6607" *)
  wire _04412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6608" *)
  wire _04413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6608" *)
  wire _04414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6609" *)
  wire _04415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6609" *)
  wire _04416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6610" *)
  wire _04417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6610" *)
  wire _04418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6611" *)
  wire _04419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6611" *)
  wire _04420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6612" *)
  wire _04421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6612" *)
  wire _04422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6613" *)
  wire _04423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6613" *)
  wire _04424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6614" *)
  wire _04425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6614" *)
  wire _04426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6615" *)
  wire _04427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6615" *)
  wire _04428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6616" *)
  wire _04429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6616" *)
  wire _04430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6617" *)
  wire _04431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6617" *)
  wire _04432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6618" *)
  wire _04433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6618" *)
  wire _04434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6619" *)
  wire _04435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6619" *)
  wire _04436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6620" *)
  wire _04437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6620" *)
  wire _04438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6621" *)
  wire _04439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6621" *)
  wire _04440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6622" *)
  wire _04441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6622" *)
  wire _04442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6623" *)
  wire _04443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6623" *)
  wire _04444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6624" *)
  wire _04445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6624" *)
  wire _04446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6625" *)
  wire _04447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6625" *)
  wire _04448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6626" *)
  wire _04449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6626" *)
  wire _04450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6627" *)
  wire _04451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6627" *)
  wire _04452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6628" *)
  wire _04453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6628" *)
  wire _04454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6629" *)
  wire _04455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6629" *)
  wire _04456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6630" *)
  wire _04457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6630" *)
  wire _04458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6631" *)
  wire _04459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6631" *)
  wire _04460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6632" *)
  wire _04461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6632" *)
  wire _04462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6633" *)
  wire _04463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6633" *)
  wire _04464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6634" *)
  wire _04465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6634" *)
  wire _04466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6635" *)
  wire _04467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6635" *)
  wire _04468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6636" *)
  wire _04469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6636" *)
  wire _04470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6637" *)
  wire _04471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6637" *)
  wire _04472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6638" *)
  wire _04473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6638" *)
  wire _04474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6639" *)
  wire _04475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6639" *)
  wire _04476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6640" *)
  wire _04477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6640" *)
  wire _04478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6641" *)
  wire _04479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6641" *)
  wire _04480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6642" *)
  wire _04481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6642" *)
  wire _04482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6643" *)
  wire _04483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6643" *)
  wire _04484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6644" *)
  wire _04485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6644" *)
  wire _04486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6645" *)
  wire _04487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6645" *)
  wire _04488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6646" *)
  wire _04489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6646" *)
  wire _04490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6647" *)
  wire _04491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6647" *)
  wire _04492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6648" *)
  wire _04493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6648" *)
  wire _04494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6649" *)
  wire _04495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6649" *)
  wire _04496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6650" *)
  wire _04497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6650" *)
  wire _04498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6651" *)
  wire _04499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6651" *)
  wire _04500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6652" *)
  wire _04501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6652" *)
  wire _04502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6653" *)
  wire _04503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6653" *)
  wire _04504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6654" *)
  wire _04505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6654" *)
  wire _04506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6655" *)
  wire _04507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6655" *)
  wire _04508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6656" *)
  wire _04509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6656" *)
  wire _04510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6657" *)
  wire _04511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6657" *)
  wire _04512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6658" *)
  wire _04513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6658" *)
  wire _04514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6659" *)
  wire _04515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6659" *)
  wire _04516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6660" *)
  wire _04517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6660" *)
  wire _04518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6661" *)
  wire _04519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6661" *)
  wire _04520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6662" *)
  wire _04521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6662" *)
  wire _04522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6663" *)
  wire _04523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6663" *)
  wire _04524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6664" *)
  wire _04525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6664" *)
  wire _04526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6665" *)
  wire _04527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6665" *)
  wire _04528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6666" *)
  wire _04529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6666" *)
  wire _04530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6667" *)
  wire _04531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6667" *)
  wire _04532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6668" *)
  wire _04533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6668" *)
  wire _04534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6669" *)
  wire _04535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6669" *)
  wire _04536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6670" *)
  wire _04537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6670" *)
  wire _04538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6671" *)
  wire _04539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6671" *)
  wire _04540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6672" *)
  wire _04541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6672" *)
  wire _04542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6673" *)
  wire _04543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6673" *)
  wire _04544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6674" *)
  wire _04545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6674" *)
  wire _04546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6675" *)
  wire _04547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6675" *)
  wire _04548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6676" *)
  wire _04549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6676" *)
  wire _04550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6677" *)
  wire _04551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6677" *)
  wire _04552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6678" *)
  wire _04553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6678" *)
  wire _04554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6679" *)
  wire _04555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6679" *)
  wire _04556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6680" *)
  wire _04557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6680" *)
  wire _04558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6681" *)
  wire _04559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6681" *)
  wire _04560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6682" *)
  wire _04561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6682" *)
  wire _04562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6683" *)
  wire _04563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6683" *)
  wire _04564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6684" *)
  wire _04565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6684" *)
  wire _04566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6685" *)
  wire _04567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6685" *)
  wire _04568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6686" *)
  wire _04569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6686" *)
  wire _04570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6687" *)
  wire _04571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6687" *)
  wire _04572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6688" *)
  wire _04573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6688" *)
  wire _04574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6689" *)
  wire _04575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6689" *)
  wire _04576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6690" *)
  wire _04577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6690" *)
  wire _04578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6691" *)
  wire _04579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6691" *)
  wire _04580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6692" *)
  wire _04581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6692" *)
  wire _04582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6693" *)
  wire _04583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6693" *)
  wire _04584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6694" *)
  wire _04585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6694" *)
  wire _04586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6695" *)
  wire _04587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6695" *)
  wire _04588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6696" *)
  wire _04589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6696" *)
  wire _04590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6697" *)
  wire _04591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6697" *)
  wire _04592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6698" *)
  wire _04593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6698" *)
  wire _04594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6699" *)
  wire _04595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6699" *)
  wire _04596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6700" *)
  wire _04597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6700" *)
  wire _04598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6701" *)
  wire _04599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6701" *)
  wire _04600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6702" *)
  wire _04601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6702" *)
  wire _04602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6703" *)
  wire _04603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6703" *)
  wire _04604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6704" *)
  wire _04605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6704" *)
  wire _04606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6705" *)
  wire _04607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6705" *)
  wire _04608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6706" *)
  wire _04609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6706" *)
  wire _04610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6707" *)
  wire _04611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6707" *)
  wire _04612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6708" *)
  wire _04613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6708" *)
  wire _04614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6709" *)
  wire _04615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6709" *)
  wire _04616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6710" *)
  wire _04617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6710" *)
  wire _04618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6711" *)
  wire _04619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6711" *)
  wire _04620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6712" *)
  wire _04621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6712" *)
  wire _04622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6713" *)
  wire _04623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6713" *)
  wire _04624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6714" *)
  wire _04625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6714" *)
  wire _04626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6715" *)
  wire _04627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6715" *)
  wire _04628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6716" *)
  wire _04629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6716" *)
  wire _04630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6717" *)
  wire _04631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6717" *)
  wire _04632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6718" *)
  wire _04633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6718" *)
  wire _04634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6719" *)
  wire _04635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6719" *)
  wire _04636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6720" *)
  wire _04637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6720" *)
  wire _04638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6721" *)
  wire _04639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6721" *)
  wire _04640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6722" *)
  wire _04641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6722" *)
  wire _04642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6723" *)
  wire _04643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6723" *)
  wire _04644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6724" *)
  wire _04645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6724" *)
  wire _04646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6725" *)
  wire _04647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6725" *)
  wire _04648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6726" *)
  wire _04649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6726" *)
  wire _04650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6727" *)
  wire _04651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6727" *)
  wire _04652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6728" *)
  wire _04653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6728" *)
  wire _04654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6729" *)
  wire _04655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6729" *)
  wire _04656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6730" *)
  wire _04657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6730" *)
  wire _04658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6731" *)
  wire _04659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6731" *)
  wire _04660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6732" *)
  wire _04661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6732" *)
  wire _04662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6733" *)
  wire _04663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6733" *)
  wire _04664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6734" *)
  wire _04665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6734" *)
  wire _04666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6735" *)
  wire _04667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6735" *)
  wire _04668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6736" *)
  wire _04669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6736" *)
  wire _04670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6737" *)
  wire _04671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6737" *)
  wire _04672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6738" *)
  wire _04673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6738" *)
  wire _04674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6739" *)
  wire _04675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6739" *)
  wire _04676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6740" *)
  wire _04677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6740" *)
  wire _04678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6741" *)
  wire _04679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6741" *)
  wire _04680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6742" *)
  wire _04681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6742" *)
  wire _04682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6743" *)
  wire _04683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6743" *)
  wire _04684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6744" *)
  wire _04685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6744" *)
  wire _04686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6745" *)
  wire _04687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6745" *)
  wire _04688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6746" *)
  wire _04689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6746" *)
  wire _04690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6747" *)
  wire _04691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6747" *)
  wire _04692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6748" *)
  wire _04693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6748" *)
  wire _04694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6749" *)
  wire _04695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6749" *)
  wire _04696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6750" *)
  wire _04697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6750" *)
  wire _04698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6751" *)
  wire _04699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6751" *)
  wire _04700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6752" *)
  wire _04701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6752" *)
  wire _04702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6753" *)
  wire _04703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6753" *)
  wire _04704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6754" *)
  wire _04705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6754" *)
  wire _04706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6755" *)
  wire _04707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6755" *)
  wire _04708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6756" *)
  wire _04709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6756" *)
  wire _04710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6757" *)
  wire _04711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6757" *)
  wire _04712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6758" *)
  wire _04713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6758" *)
  wire _04714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6759" *)
  wire _04715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6759" *)
  wire _04716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6760" *)
  wire _04717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6760" *)
  wire _04718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6761" *)
  wire _04719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6761" *)
  wire _04720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6762" *)
  wire _04721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6762" *)
  wire _04722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6763" *)
  wire _04723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6763" *)
  wire _04724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6764" *)
  wire _04725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6764" *)
  wire _04726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6765" *)
  wire _04727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6765" *)
  wire _04728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6766" *)
  wire _04729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6766" *)
  wire _04730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6767" *)
  wire _04731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6767" *)
  wire _04732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6768" *)
  wire _04733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6768" *)
  wire _04734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6769" *)
  wire _04735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6769" *)
  wire _04736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6770" *)
  wire _04737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6770" *)
  wire _04738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6771" *)
  wire _04739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6771" *)
  wire _04740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6772" *)
  wire _04741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6772" *)
  wire _04742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6773" *)
  wire _04743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6773" *)
  wire _04744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6774" *)
  wire _04745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6774" *)
  wire _04746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6775" *)
  wire _04747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6775" *)
  wire _04748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6776" *)
  wire _04749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6776" *)
  wire _04750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6777" *)
  wire _04751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6777" *)
  wire _04752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6778" *)
  wire _04753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6778" *)
  wire _04754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6779" *)
  wire _04755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6779" *)
  wire _04756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6780" *)
  wire _04757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6780" *)
  wire _04758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6781" *)
  wire _04759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6781" *)
  wire _04760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6782" *)
  wire _04761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6782" *)
  wire _04762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6783" *)
  wire _04763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6783" *)
  wire _04764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6784" *)
  wire _04765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6784" *)
  wire _04766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6785" *)
  wire _04767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6785" *)
  wire _04768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6786" *)
  wire _04769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6786" *)
  wire _04770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6787" *)
  wire _04771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6787" *)
  wire _04772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6788" *)
  wire _04773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6788" *)
  wire _04774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6789" *)
  wire _04775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6789" *)
  wire _04776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6790" *)
  wire _04777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6790" *)
  wire _04778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6791" *)
  wire _04779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6791" *)
  wire _04780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6792" *)
  wire _04781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6792" *)
  wire _04782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6793" *)
  wire _04783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6793" *)
  wire _04784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6794" *)
  wire _04785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6794" *)
  wire _04786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6795" *)
  wire _04787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6795" *)
  wire _04788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6796" *)
  wire _04789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6796" *)
  wire _04790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6797" *)
  wire _04791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6797" *)
  wire _04792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6798" *)
  wire _04793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6798" *)
  wire _04794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6799" *)
  wire _04795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6799" *)
  wire _04796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6800" *)
  wire _04797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6800" *)
  wire _04798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6801" *)
  wire _04799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6801" *)
  wire _04800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6802" *)
  wire _04801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6802" *)
  wire _04802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6803" *)
  wire _04803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6803" *)
  wire _04804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6804" *)
  wire _04805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6804" *)
  wire _04806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6805" *)
  wire _04807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6805" *)
  wire _04808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6806" *)
  wire _04809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6806" *)
  wire _04810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6807" *)
  wire _04811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6807" *)
  wire _04812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6808" *)
  wire _04813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6808" *)
  wire _04814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6809" *)
  wire _04815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6809" *)
  wire _04816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6810" *)
  wire _04817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6810" *)
  wire _04818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6811" *)
  wire _04819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6811" *)
  wire _04820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6812" *)
  wire _04821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6812" *)
  wire _04822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6813" *)
  wire _04823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6813" *)
  wire _04824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6814" *)
  wire _04825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6814" *)
  wire _04826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6815" *)
  wire _04827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6815" *)
  wire _04828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6816" *)
  wire _04829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6816" *)
  wire _04830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6817" *)
  wire _04831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6817" *)
  wire _04832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6818" *)
  wire _04833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6818" *)
  wire _04834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6819" *)
  wire _04835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6819" *)
  wire _04836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6820" *)
  wire _04837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6820" *)
  wire _04838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6821" *)
  wire _04839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6821" *)
  wire _04840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6822" *)
  wire _04841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6822" *)
  wire _04842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6823" *)
  wire _04843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6823" *)
  wire _04844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6824" *)
  wire _04845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6824" *)
  wire _04846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6825" *)
  wire _04847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6825" *)
  wire _04848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6826" *)
  wire _04849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6826" *)
  wire _04850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6827" *)
  wire _04851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6827" *)
  wire _04852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6828" *)
  wire _04853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6828" *)
  wire _04854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6829" *)
  wire _04855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6829" *)
  wire _04856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6830" *)
  wire _04857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6830" *)
  wire _04858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6831" *)
  wire _04859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6831" *)
  wire _04860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6832" *)
  wire _04861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6832" *)
  wire _04862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6833" *)
  wire _04863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6833" *)
  wire _04864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6834" *)
  wire _04865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6834" *)
  wire _04866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6835" *)
  wire _04867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6835" *)
  wire _04868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6836" *)
  wire _04869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6836" *)
  wire _04870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6837" *)
  wire _04871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6837" *)
  wire _04872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6838" *)
  wire _04873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6838" *)
  wire _04874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6839" *)
  wire _04875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6839" *)
  wire _04876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6840" *)
  wire _04877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6840" *)
  wire _04878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6841" *)
  wire _04879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6841" *)
  wire _04880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6842" *)
  wire _04881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6842" *)
  wire _04882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6843" *)
  wire _04883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6843" *)
  wire _04884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6844" *)
  wire _04885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6844" *)
  wire _04886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6845" *)
  wire _04887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6845" *)
  wire _04888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6846" *)
  wire _04889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6846" *)
  wire _04890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6847" *)
  wire _04891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6847" *)
  wire _04892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6848" *)
  wire _04893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6848" *)
  wire _04894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6849" *)
  wire _04895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6849" *)
  wire _04896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6850" *)
  wire _04897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6850" *)
  wire _04898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6851" *)
  wire _04899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6851" *)
  wire _04900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6852" *)
  wire _04901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6852" *)
  wire _04902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6853" *)
  wire _04903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6853" *)
  wire _04904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6854" *)
  wire _04905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6854" *)
  wire _04906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6855" *)
  wire _04907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6855" *)
  wire _04908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6856" *)
  wire _04909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6856" *)
  wire _04910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6857" *)
  wire _04911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6857" *)
  wire _04912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6858" *)
  wire _04913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6858" *)
  wire _04914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6859" *)
  wire _04915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6859" *)
  wire _04916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6860" *)
  wire _04917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6860" *)
  wire _04918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6861" *)
  wire _04919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6861" *)
  wire _04920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6862" *)
  wire _04921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6862" *)
  wire _04922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6863" *)
  wire _04923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6863" *)
  wire _04924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6864" *)
  wire _04925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6864" *)
  wire _04926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6865" *)
  wire _04927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6865" *)
  wire _04928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6866" *)
  wire _04929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6866" *)
  wire _04930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6867" *)
  wire _04931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6867" *)
  wire _04932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6868" *)
  wire _04933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6868" *)
  wire _04934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6869" *)
  wire _04935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6869" *)
  wire _04936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6870" *)
  wire _04937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6870" *)
  wire _04938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6871" *)
  wire _04939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6871" *)
  wire _04940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6872" *)
  wire _04941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6872" *)
  wire _04942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6873" *)
  wire _04943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6873" *)
  wire _04944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6874" *)
  wire _04945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6874" *)
  wire _04946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6875" *)
  wire _04947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6875" *)
  wire _04948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6876" *)
  wire _04949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6876" *)
  wire _04950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6877" *)
  wire _04951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6877" *)
  wire _04952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6878" *)
  wire _04953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6878" *)
  wire _04954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6879" *)
  wire _04955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6879" *)
  wire _04956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6880" *)
  wire _04957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6880" *)
  wire _04958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6881" *)
  wire _04959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6881" *)
  wire _04960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6882" *)
  wire _04961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6882" *)
  wire _04962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6883" *)
  wire _04963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6883" *)
  wire _04964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6884" *)
  wire _04965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6884" *)
  wire _04966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6885" *)
  wire _04967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6885" *)
  wire _04968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6886" *)
  wire _04969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6886" *)
  wire _04970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6887" *)
  wire _04971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6887" *)
  wire _04972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6888" *)
  wire _04973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6888" *)
  wire _04974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6889" *)
  wire _04975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6889" *)
  wire _04976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6890" *)
  wire _04977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6890" *)
  wire _04978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6891" *)
  wire _04979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6891" *)
  wire _04980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6892" *)
  wire _04981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6892" *)
  wire _04982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6893" *)
  wire _04983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6893" *)
  wire _04984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6894" *)
  wire _04985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6894" *)
  wire _04986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6895" *)
  wire _04987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6895" *)
  wire _04988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6896" *)
  wire _04989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6896" *)
  wire _04990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6897" *)
  wire _04991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6897" *)
  wire _04992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6898" *)
  wire _04993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6898" *)
  wire _04994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6899" *)
  wire _04995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6899" *)
  wire _04996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6900" *)
  wire _04997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6900" *)
  wire _04998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6901" *)
  wire _04999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6901" *)
  wire _05000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6902" *)
  wire _05001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6902" *)
  wire _05002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6903" *)
  wire _05003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6903" *)
  wire _05004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6904" *)
  wire _05005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6904" *)
  wire _05006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6905" *)
  wire _05007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6905" *)
  wire _05008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6906" *)
  wire _05009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6906" *)
  wire _05010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6907" *)
  wire _05011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6907" *)
  wire _05012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6908" *)
  wire _05013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6908" *)
  wire _05014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6909" *)
  wire _05015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6909" *)
  wire _05016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6910" *)
  wire _05017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6910" *)
  wire _05018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6911" *)
  wire _05019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6911" *)
  wire _05020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6912" *)
  wire _05021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6912" *)
  wire _05022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6913" *)
  wire _05023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6913" *)
  wire _05024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6914" *)
  wire _05025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6914" *)
  wire _05026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6915" *)
  wire _05027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6915" *)
  wire _05028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6916" *)
  wire _05029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6916" *)
  wire _05030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6917" *)
  wire _05031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6917" *)
  wire _05032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6918" *)
  wire _05033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6918" *)
  wire _05034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6919" *)
  wire _05035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6919" *)
  wire _05036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6920" *)
  wire _05037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6920" *)
  wire _05038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6921" *)
  wire _05039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6921" *)
  wire _05040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6922" *)
  wire _05041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6922" *)
  wire _05042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6923" *)
  wire _05043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6923" *)
  wire _05044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6924" *)
  wire _05045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6924" *)
  wire _05046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6925" *)
  wire _05047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6925" *)
  wire _05048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6926" *)
  wire _05049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6926" *)
  wire _05050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6927" *)
  wire _05051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6927" *)
  wire _05052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6928" *)
  wire _05053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6928" *)
  wire _05054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6929" *)
  wire _05055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6929" *)
  wire _05056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6930" *)
  wire _05057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6930" *)
  wire _05058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6931" *)
  wire _05059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6931" *)
  wire _05060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6932" *)
  wire _05061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6932" *)
  wire _05062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6933" *)
  wire _05063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6933" *)
  wire _05064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6934" *)
  wire _05065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6934" *)
  wire _05066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6935" *)
  wire _05067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6935" *)
  wire _05068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6936" *)
  wire _05069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6936" *)
  wire _05070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6937" *)
  wire _05071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6937" *)
  wire _05072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6938" *)
  wire _05073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6938" *)
  wire _05074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6939" *)
  wire _05075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6939" *)
  wire _05076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6940" *)
  wire _05077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6940" *)
  wire _05078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6941" *)
  wire _05079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6941" *)
  wire _05080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6942" *)
  wire _05081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6942" *)
  wire _05082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6943" *)
  wire _05083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6943" *)
  wire _05084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6944" *)
  wire _05085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6944" *)
  wire _05086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6945" *)
  wire _05087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6945" *)
  wire _05088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6946" *)
  wire _05089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6946" *)
  wire _05090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6947" *)
  wire _05091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6947" *)
  wire _05092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6948" *)
  wire _05093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6948" *)
  wire _05094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6949" *)
  wire _05095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6949" *)
  wire _05096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6950" *)
  wire _05097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6950" *)
  wire _05098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6951" *)
  wire _05099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6951" *)
  wire _05100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6952" *)
  wire _05101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6952" *)
  wire _05102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6953" *)
  wire _05103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6953" *)
  wire _05104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6954" *)
  wire _05105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6954" *)
  wire _05106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6955" *)
  wire _05107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6955" *)
  wire _05108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6956" *)
  wire _05109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6956" *)
  wire _05110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6957" *)
  wire _05111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6957" *)
  wire _05112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6958" *)
  wire _05113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6958" *)
  wire _05114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6959" *)
  wire _05115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6959" *)
  wire _05116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6960" *)
  wire _05117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6960" *)
  wire _05118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6961" *)
  wire _05119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6961" *)
  wire _05120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6962" *)
  wire _05121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6962" *)
  wire _05122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6963" *)
  wire _05123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6963" *)
  wire _05124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6964" *)
  wire _05125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6964" *)
  wire _05126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6965" *)
  wire _05127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6965" *)
  wire _05128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6966" *)
  wire _05129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6966" *)
  wire _05130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6967" *)
  wire _05131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6967" *)
  wire _05132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6968" *)
  wire _05133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6968" *)
  wire _05134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6969" *)
  wire _05135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6969" *)
  wire _05136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6970" *)
  wire _05137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6970" *)
  wire _05138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6971" *)
  wire _05139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6971" *)
  wire _05140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6972" *)
  wire _05141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6972" *)
  wire _05142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6973" *)
  wire _05143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6973" *)
  wire _05144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6974" *)
  wire _05145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6974" *)
  wire _05146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6975" *)
  wire _05147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6975" *)
  wire _05148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6976" *)
  wire _05149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6976" *)
  wire _05150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6977" *)
  wire _05151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6977" *)
  wire _05152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6978" *)
  wire _05153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6978" *)
  wire _05154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6979" *)
  wire _05155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6979" *)
  wire _05156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6980" *)
  wire _05157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6980" *)
  wire _05158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6981" *)
  wire _05159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6981" *)
  wire _05160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6982" *)
  wire _05161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6982" *)
  wire _05162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6983" *)
  wire _05163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6983" *)
  wire _05164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6984" *)
  wire _05165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6984" *)
  wire _05166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6985" *)
  wire _05167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6985" *)
  wire _05168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6986" *)
  wire _05169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6986" *)
  wire _05170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6987" *)
  wire _05171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6987" *)
  wire _05172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6988" *)
  wire _05173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6988" *)
  wire _05174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6989" *)
  wire _05175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6989" *)
  wire _05176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6990" *)
  wire _05177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6990" *)
  wire _05178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6991" *)
  wire _05179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6991" *)
  wire _05180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6992" *)
  wire _05181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6992" *)
  wire _05182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6993" *)
  wire _05183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6993" *)
  wire _05184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6994" *)
  wire _05185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6994" *)
  wire _05186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6995" *)
  wire _05187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6995" *)
  wire _05188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6996" *)
  wire _05189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6996" *)
  wire _05190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6997" *)
  wire _05191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6997" *)
  wire _05192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6998" *)
  wire _05193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6998" *)
  wire _05194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6999" *)
  wire _05195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6999" *)
  wire _05196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7000" *)
  wire _05197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7000" *)
  wire _05198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7001" *)
  wire _05199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7001" *)
  wire _05200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7002" *)
  wire _05201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7002" *)
  wire _05202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7003" *)
  wire _05203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7003" *)
  wire _05204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7004" *)
  wire _05205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7004" *)
  wire _05206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7005" *)
  wire _05207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7005" *)
  wire _05208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7006" *)
  wire _05209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7006" *)
  wire _05210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7007" *)
  wire _05211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7007" *)
  wire _05212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7008" *)
  wire _05213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7008" *)
  wire _05214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7009" *)
  wire _05215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7009" *)
  wire _05216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7010" *)
  wire _05217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7010" *)
  wire _05218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7011" *)
  wire _05219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7011" *)
  wire _05220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7012" *)
  wire _05221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7012" *)
  wire _05222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7013" *)
  wire _05223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7013" *)
  wire _05224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7014" *)
  wire _05225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7014" *)
  wire _05226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7015" *)
  wire _05227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7015" *)
  wire _05228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7016" *)
  wire _05229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7016" *)
  wire _05230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7017" *)
  wire _05231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7017" *)
  wire _05232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7018" *)
  wire _05233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7018" *)
  wire _05234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7019" *)
  wire _05235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7019" *)
  wire _05236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7020" *)
  wire _05237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7020" *)
  wire _05238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7021" *)
  wire _05239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7021" *)
  wire _05240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7022" *)
  wire _05241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7022" *)
  wire _05242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7023" *)
  wire _05243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7023" *)
  wire _05244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7024" *)
  wire _05245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7024" *)
  wire _05246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7025" *)
  wire _05247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7025" *)
  wire _05248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7026" *)
  wire _05249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7026" *)
  wire _05250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7027" *)
  wire _05251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7027" *)
  wire _05252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7028" *)
  wire _05253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7028" *)
  wire _05254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7029" *)
  wire _05255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7029" *)
  wire _05256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7030" *)
  wire _05257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7030" *)
  wire _05258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7031" *)
  wire _05259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7031" *)
  wire _05260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7032" *)
  wire _05261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7032" *)
  wire _05262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7033" *)
  wire _05263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7033" *)
  wire _05264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7034" *)
  wire _05265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7034" *)
  wire _05266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7035" *)
  wire _05267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7035" *)
  wire _05268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7036" *)
  wire _05269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7036" *)
  wire _05270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7037" *)
  wire _05271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7037" *)
  wire _05272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7038" *)
  wire _05273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7038" *)
  wire _05274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7039" *)
  wire _05275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7039" *)
  wire _05276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7040" *)
  wire _05277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7040" *)
  wire _05278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7041" *)
  wire _05279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7041" *)
  wire _05280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7042" *)
  wire _05281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7042" *)
  wire _05282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7043" *)
  wire _05283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7043" *)
  wire _05284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7044" *)
  wire _05285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7044" *)
  wire _05286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7045" *)
  wire _05287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7045" *)
  wire _05288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7046" *)
  wire _05289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7046" *)
  wire _05290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7112" *)
  wire _05291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7112" *)
  wire _05292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7114" *)
  wire _05293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7116" *)
  wire _05294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7117" *)
  wire _05295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7117" *)
  wire _05296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7117" *)
  wire _05297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7117" *)
  wire _05298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7120" *)
  wire _05299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7120" *)
  wire _05300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7120" *)
  wire _05301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7123" *)
  wire _05302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7124" *)
  wire _05303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7127" *)
  wire _05304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7127" *)
  wire _05305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7129" *)
  wire _05306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7131" *)
  wire _05307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7132" *)
  wire _05308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7132" *)
  wire _05309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7132" *)
  wire _05310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7132" *)
  wire _05311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7135" *)
  wire _05312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7135" *)
  wire _05313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7135" *)
  wire _05314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7138" *)
  wire _05315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7139" *)
  wire _05316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7142" *)
  wire _05317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7142" *)
  wire _05318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7144" *)
  wire _05319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7146" *)
  wire _05320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7147" *)
  wire _05321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7147" *)
  wire _05322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7147" *)
  wire _05323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7147" *)
  wire _05324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7150" *)
  wire _05325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7150" *)
  wire _05326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7150" *)
  wire _05327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7153" *)
  wire _05328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7154" *)
  wire _05329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7156" *)
  wire _05330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7156" *)
  wire _05331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7157" *)
  wire _05332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7157" *)
  wire _05333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7157" *)
  wire _05334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7159" *)
  wire _05335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7159" *)
  wire _05336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7162" *)
  wire _05337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7163" *)
  wire _05338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7163" *)
  wire _05339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7163" *)
  wire _05340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7163" *)
  wire _05341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7167" *)
  wire _05342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7167" *)
  wire _05343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7170" *)
  wire _05344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7171" *)
  wire _05345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7177" *)
  wire _05346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7184" *)
  wire _05347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7184" *)
  wire _05348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7185" *)
  wire _05349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7190" *)
  wire _05350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7190" *)
  wire _05351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7190" *)
  wire _05352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7194" *)
  wire _05353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7194" *)
  wire _05354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7195" *)
  wire _05355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7195" *)
  wire _05356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7196" *)
  wire _05357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7197" *)
  wire _05358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7197" *)
  wire _05359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7199" *)
  wire _05360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7199" *)
  wire _05361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7206" *)
  wire _05362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7206" *)
  wire _05363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7207" *)
  wire _05364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7207" *)
  wire _05365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7209" *)
  wire _05366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7209" *)
  wire _05367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7209" *)
  wire _05368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7212" *)
  wire _05369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7212" *)
  wire _05370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7215" *)
  wire _05371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7215" *)
  wire _05372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7218" *)
  wire _05373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7218" *)
  wire _05374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7218" *)
  wire _05375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7221" *)
  wire _05376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7222" *)
  wire _05377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7222" *)
  wire _05378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7223" *)
  wire _05379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7224" *)
  wire _05380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7224" *)
  wire _05381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7226" *)
  wire _05382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7226" *)
  wire _05383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7228" *)
  wire _05384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7233" *)
  wire _05385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7233" *)
  wire _05386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7234" *)
  wire _05387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7234" *)
  wire _05388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7236" *)
  wire _05389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7236" *)
  wire _05390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7236" *)
  wire _05391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7240" *)
  wire _05392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7240" *)
  wire _05393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7243" *)
  wire _05394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7243" *)
  wire _05395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7246" *)
  wire _05396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7246" *)
  wire _05397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7246" *)
  wire _05398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7249" *)
  wire _05399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7250" *)
  wire _05400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7250" *)
  wire _05401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7251" *)
  wire _05402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7252" *)
  wire _05403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7252" *)
  wire _05404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7254" *)
  wire _05405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7254" *)
  wire _05406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7256" *)
  wire _05407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7261" *)
  wire _05408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7261" *)
  wire _05409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7262" *)
  wire _05410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7262" *)
  wire _05411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7264" *)
  wire _05412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7264" *)
  wire _05413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7264" *)
  wire _05414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7268" *)
  wire _05415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7268" *)
  wire _05416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7273" *)
  wire _05417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7273" *)
  wire _05418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7274" *)
  wire _05419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7275" *)
  wire _05420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7277" *)
  wire _05421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7277" *)
  wire _05422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7277" *)
  wire _05423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7281" *)
  wire _05424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7282" *)
  wire _05425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7282" *)
  wire _05426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7282" *)
  wire _05427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7284" *)
  wire _05428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7284" *)
  wire _05429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7284" *)
  wire _05430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7286" *)
  wire _05431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7290" *)
  wire _05432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7291" *)
  wire _05433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7291" *)
  wire _05434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7293" *)
  wire _05435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7293" *)
  wire _05436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7293" *)
  wire _05437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7296" *)
  wire _05438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7296" *)
  wire _05439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7296" *)
  wire _05440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7296" *)
  wire _05441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7337" *)
  wire _05442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7338" *)
  wire _05443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7339" *)
  wire _05444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7342" *)
  wire _05445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7343" *)
  wire _05446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7344" *)
  wire _05447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7345" *)
  wire _05448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7346" *)
  wire _05449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7347" *)
  wire _05450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7348" *)
  wire _05451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7349" *)
  wire _05452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7350" *)
  wire _05453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7351" *)
  wire _05454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7351" *)
  wire _05455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7352" *)
  wire _05456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7353" *)
  wire _05457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7354" *)
  wire _05458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7360" *)
  wire _05459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7361" *)
  wire _05460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7362" *)
  wire _05461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7363" *)
  wire _05462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7370" *)
  wire _05463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7473" *)
  wire _05464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7481" *)
  wire _05465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7489" *)
  wire _05466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7745" *)
  wire _05467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8382" *)
  wire _05468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8430" *)
  wire _05469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8497" *)
  wire _05470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8539" *)
  wire _05471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8605" *)
  wire _05472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8605" *)
  wire _05473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8670" *)
  wire _05474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8670" *)
  wire _05475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8735" *)
  wire _05476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8735" *)
  wire _05477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8776" *)
  wire _05478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8776" *)
  wire _05479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8784" *)
  wire _05480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8784" *)
  wire _05481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8804" *)
  wire _05482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8804" *)
  wire _05483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8812" *)
  wire _05484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8812" *)
  wire _05485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8832" *)
  wire _05486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8832" *)
  wire _05487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8840" *)
  wire _05488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8840" *)
  wire _05489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8860" *)
  wire _05490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8860" *)
  wire _05491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8868" *)
  wire _05492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8868" *)
  wire _05493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8879" *)
  wire _05494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8880" *)
  wire _05495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8880" *)
  wire _05496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8890" *)
  wire _05497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8902" *)
  wire _05498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8911" *)
  wire _05499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8911" *)
  wire _05500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8921" *)
  wire _05501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8932" *)
  wire _05502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8932" *)
  wire _05503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8942" *)
  wire _05504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8954" *)
  wire _05505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8954" *)
  wire _05506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8964" *)
  wire _05507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8983" *)
  wire _05508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8999" *)
  wire _05509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9015" *)
  wire _05510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9031" *)
  wire _05511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9079" *)
  wire _05512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *)
  wire _05513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *)
  wire _05514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *)
  wire _05515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *)
  wire _05516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *)
  wire _05517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9097" *)
  wire _05518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9098" *)
  wire _05519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9098" *)
  wire _05520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *)
  wire _05521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *)
  wire _05522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *)
  wire _05523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *)
  wire _05524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *)
  wire _05525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9116" *)
  wire _05526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9117" *)
  wire _05527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9117" *)
  wire _05528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *)
  wire _05529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *)
  wire _05530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *)
  wire _05531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *)
  wire _05532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *)
  wire _05533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9135" *)
  wire _05534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9136" *)
  wire _05535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9136" *)
  wire _05536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9145" *)
  wire _05537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9145" *)
  wire _05538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9146" *)
  wire _05539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9146" *)
  wire _05540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9146" *)
  wire _05541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9154" *)
  wire _05542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9155" *)
  wire _05543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9155" *)
  wire _05544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9161" *)
  wire _05545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9161" *)
  wire _05546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9169" *)
  wire _05547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9169" *)
  wire _05548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9176" *)
  wire _05549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9176" *)
  wire _05550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9184" *)
  wire _05551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9184" *)
  wire _05552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9191" *)
  wire _05553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9191" *)
  wire _05554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9199" *)
  wire _05555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9199" *)
  wire _05556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9205" *)
  wire _05557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9206" *)
  wire _05558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9213" *)
  wire _05559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9214" *)
  wire _05560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9224" *)
  wire _05561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9242" *)
  wire _05562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9260" *)
  wire _05563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9278" *)
  wire _05564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9292" *)
  wire _05565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9295" *)
  wire _05566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9295" *)
  wire _05567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9295" *)
  wire _05568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9296" *)
  wire _05569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9299" *)
  wire _05570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9302" *)
  wire _05571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9302" *)
  wire _05572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9303" *)
  wire _05573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9306" *)
  wire _05574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9309" *)
  wire _05575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9309" *)
  wire _05576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9310" *)
  wire _05577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9313" *)
  wire _05578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9316" *)
  wire _05579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9316" *)
  wire _05580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9316" *)
  wire _05581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9317" *)
  wire _05582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9320" *)
  wire _05583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9320" *)
  wire _05584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9320" *)
  wire _05585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9321" *)
  wire _05586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9322" *)
  wire _05587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9324" *)
  wire _05588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9324" *)
  wire _05589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9327" *)
  wire _05590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9328" *)
  wire _05591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9331" *)
  wire _05592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9335" *)
  wire _05593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9340" *)
  wire _05594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9347" *)
  wire _05595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9350" *)
  wire _05596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9350" *)
  wire _05597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9350" *)
  wire _05598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9350" *)
  wire _05599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9352" *)
  wire _05600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9352" *)
  wire _05601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9353" *)
  wire _05602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9353" *)
  wire _05603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9356" *)
  wire _05604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9356" *)
  wire _05605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9357" *)
  wire _05606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9359" *)
  wire _05607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9360" *)
  wire _05608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9362" *)
  wire _05609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9362" *)
  wire _05610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9365" *)
  wire _05611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9366" *)
  wire _05612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9371" *)
  wire _05613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9374" *)
  wire _05614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9375" *)
  wire _05615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9375" *)
  wire _05616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9378" *)
  wire _05617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9380" *)
  wire _05618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9383" *)
  wire _05619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9383" *)
  wire _05620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9383" *)
  wire _05621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9384" *)
  wire _05622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9388" *)
  wire _05623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9388" *)
  wire _05624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9390" *)
  wire _05625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9390" *)
  wire _05626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9395" *)
  wire _05627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9400" *)
  wire _05628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *)
  wire _05629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *)
  wire _05630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *)
  wire _05631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *)
  wire _05632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9405" *)
  wire _05633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9406" *)
  wire _05634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9406" *)
  wire _05635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9406" *)
  wire _05636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9407" *)
  wire _05637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9407" *)
  wire _05638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9407" *)
  wire _05639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9409" *)
  wire _05640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9409" *)
  wire _05641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9409" *)
  wire _05642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9410" *)
  wire _05643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9410" *)
  wire _05644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9410" *)
  wire _05645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9410" *)
  wire _05646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9415" *)
  wire _05647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9415" *)
  wire _05648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9415" *)
  wire _05649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9416" *)
  wire _05650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9416" *)
  wire _05651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9416" *)
  wire _05652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9416" *)
  wire _05653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9418" *)
  wire _05654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9419" *)
  wire _05655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9419" *)
  wire _05656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9419" *)
  wire _05657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9420" *)
  wire _05658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9420" *)
  wire _05659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9420" *)
  wire _05660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9420" *)
  wire _05661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9423" *)
  wire _05662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9424" *)
  wire _05663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9425" *)
  wire _05664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9425" *)
  wire _05665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9427" *)
  wire _05666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9428" *)
  wire _05667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9428" *)
  wire _05668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9431" *)
  wire _05669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9432" *)
  wire _05670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9432" *)
  wire _05671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9435" *)
  wire _05672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9440" *)
  wire _05673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9441" *)
  wire _05674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9446" *)
  wire _05675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9451" *)
  wire _05676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9454" *)
  wire _05677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9454" *)
  wire _05678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9454" *)
  wire _05679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9454" *)
  wire _05680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9456" *)
  wire _05681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9456" *)
  wire _05682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9457" *)
  wire _05683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9457" *)
  wire _05684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9460" *)
  wire _05685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9460" *)
  wire _05686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9461" *)
  wire _05687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9463" *)
  wire _05688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9464" *)
  wire _05689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9466" *)
  wire _05690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9466" *)
  wire _05691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9469" *)
  wire _05692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9470" *)
  wire _05693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9475" *)
  wire _05694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9477" *)
  wire _05695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9477" *)
  wire _05696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9478" *)
  wire _05697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9478" *)
  wire _05698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9478" *)
  wire _05699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9479" *)
  wire _05700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9479" *)
  wire _05701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9479" *)
  wire _05702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9482" *)
  wire _05703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9484" *)
  wire _05704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9490" *)
  wire _05705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9490" *)
  wire _05706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9491" *)
  wire _05707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9492" *)
  wire _05708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9492" *)
  wire _05709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9494" *)
  wire _05710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9494" *)
  wire _05711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9494" *)
  wire _05712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9499" *)
  wire _05713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9499" *)
  wire _05714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9501" *)
  wire _05715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9507" *)
  wire _05716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9507" *)
  wire _05717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9508" *)
  wire _05718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9508" *)
  wire _05719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9511" *)
  wire _05720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9511" *)
  wire _05721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9511" *)
  wire _05722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9512" *)
  wire _05723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9512" *)
  wire _05724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9512" *)
  wire _05725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9514" *)
  wire _05726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9514" *)
  wire _05727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9515" *)
  wire _05728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9515" *)
  wire _05729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9515" *)
  wire _05730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9515" *)
  wire _05731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9520" *)
  wire _05732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9520" *)
  wire _05733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9521" *)
  wire _05734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9521" *)
  wire _05735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9521" *)
  wire _05736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9521" *)
  wire _05737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9523" *)
  wire _05738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9524" *)
  wire _05739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9524" *)
  wire _05740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9524" *)
  wire _05741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9525" *)
  wire _05742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9525" *)
  wire _05743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9525" *)
  wire _05744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9525" *)
  wire _05745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9528" *)
  wire _05746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9529" *)
  wire _05747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9530" *)
  wire _05748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9530" *)
  wire _05749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9532" *)
  wire _05750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9533" *)
  wire _05751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9533" *)
  wire _05752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9536" *)
  wire _05753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9537" *)
  wire _05754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9537" *)
  wire _05755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9540" *)
  wire _05756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9545" *)
  wire _05757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9546" *)
  wire _05758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9551" *)
  wire _05759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9556" *)
  wire _05760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9559" *)
  wire _05761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9559" *)
  wire _05762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9559" *)
  wire _05763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9559" *)
  wire _05764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9561" *)
  wire _05765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9561" *)
  wire _05766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9562" *)
  wire _05767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9562" *)
  wire _05768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9565" *)
  wire _05769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9565" *)
  wire _05770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9566" *)
  wire _05771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9568" *)
  wire _05772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9569" *)
  wire _05773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9571" *)
  wire _05774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9571" *)
  wire _05775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9574" *)
  wire _05776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9575" *)
  wire _05777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9580" *)
  wire _05778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9582" *)
  wire _05779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9582" *)
  wire _05780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9583" *)
  wire _05781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9583" *)
  wire _05782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9583" *)
  wire _05783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9584" *)
  wire _05784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9584" *)
  wire _05785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9584" *)
  wire _05786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9587" *)
  wire _05787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9589" *)
  wire _05788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9595" *)
  wire _05789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9595" *)
  wire _05790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9596" *)
  wire _05791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9597" *)
  wire _05792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9597" *)
  wire _05793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9599" *)
  wire _05794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9599" *)
  wire _05795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9599" *)
  wire _05796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9604" *)
  wire _05797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9604" *)
  wire _05798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9606" *)
  wire _05799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9612" *)
  wire _05800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9612" *)
  wire _05801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9613" *)
  wire _05802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9613" *)
  wire _05803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9616" *)
  wire _05804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9616" *)
  wire _05805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9616" *)
  wire _05806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9617" *)
  wire _05807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9617" *)
  wire _05808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9617" *)
  wire _05809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9619" *)
  wire _05810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9619" *)
  wire _05811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9620" *)
  wire _05812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9620" *)
  wire _05813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9620" *)
  wire _05814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9620" *)
  wire _05815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9625" *)
  wire _05816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9625" *)
  wire _05817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9626" *)
  wire _05818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9626" *)
  wire _05819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9626" *)
  wire _05820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9626" *)
  wire _05821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9628" *)
  wire _05822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9629" *)
  wire _05823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9629" *)
  wire _05824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9629" *)
  wire _05825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9630" *)
  wire _05826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9630" *)
  wire _05827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9630" *)
  wire _05828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9630" *)
  wire _05829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9633" *)
  wire _05830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9634" *)
  wire _05831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9635" *)
  wire _05832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9635" *)
  wire _05833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9637" *)
  wire _05834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9638" *)
  wire _05835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9638" *)
  wire _05836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9641" *)
  wire _05837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9642" *)
  wire _05838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9642" *)
  wire _05839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9645" *)
  wire _05840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9650" *)
  wire _05841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9656" *)
  wire _05842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9661" *)
  wire _05843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9664" *)
  wire _05844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9664" *)
  wire _05845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9664" *)
  wire _05846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9664" *)
  wire _05847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9666" *)
  wire _05848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9666" *)
  wire _05849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9667" *)
  wire _05850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9667" *)
  wire _05851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9670" *)
  wire _05852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9670" *)
  wire _05853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9671" *)
  wire _05854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9673" *)
  wire _05855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9674" *)
  wire _05856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9676" *)
  wire _05857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9676" *)
  wire _05858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9679" *)
  wire _05859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9680" *)
  wire _05860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9685" *)
  wire _05861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9687" *)
  wire _05862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9687" *)
  wire _05863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9688" *)
  wire _05864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9688" *)
  wire _05865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9688" *)
  wire _05866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9689" *)
  wire _05867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9689" *)
  wire _05868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9689" *)
  wire _05869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9701" *)
  wire _05870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9701" *)
  wire _05871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9702" *)
  wire _05872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9703" *)
  wire _05873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9703" *)
  wire _05874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9705" *)
  wire _05875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9705" *)
  wire _05876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9705" *)
  wire _05877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9710" *)
  wire _05878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9710" *)
  wire _05879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9712" *)
  wire _05880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9718" *)
  wire _05881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9718" *)
  wire _05882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9719" *)
  wire _05883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9719" *)
  wire _05884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9722" *)
  wire _05885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9722" *)
  wire _05886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9722" *)
  wire _05887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9723" *)
  wire _05888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9723" *)
  wire _05889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9723" *)
  wire _05890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9725" *)
  wire _05891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9725" *)
  wire _05892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9726" *)
  wire _05893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9726" *)
  wire _05894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9726" *)
  wire _05895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9726" *)
  wire _05896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9731" *)
  wire _05897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9731" *)
  wire _05898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9732" *)
  wire _05899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9732" *)
  wire _05900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9732" *)
  wire _05901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9732" *)
  wire _05902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9734" *)
  wire _05903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9735" *)
  wire _05904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9735" *)
  wire _05905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9735" *)
  wire _05906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9736" *)
  wire _05907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9736" *)
  wire _05908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9736" *)
  wire _05909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9736" *)
  wire _05910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9739" *)
  wire _05911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9741" *)
  wire _05912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9741" *)
  wire _05913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9744" *)
  wire _05914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9752" *)
  wire _05915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9753" *)
  wire _05916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9753" *)
  wire _05917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9753" *)
  wire _05918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9758" *)
  wire _05919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9758" *)
  wire _05920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9761" *)
  wire _05921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9761" *)
  wire _05922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9761" *)
  wire _05923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9771" *)
  wire _05924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9771" *)
  wire _05925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9776" *)
  wire _05926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9776" *)
  wire _05927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9779" *)
  wire _05928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9779" *)
  wire _05929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9779" *)
  wire _05930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9789" *)
  wire _05931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9789" *)
  wire _05932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9794" *)
  wire _05933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9797" *)
  wire _05934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9797" *)
  wire _05935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9801" *)
  wire _05936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9812" *)
  wire _05937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9812" *)
  wire _05938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9814" *)
  wire _05939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9814" *)
  wire _05940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9815" *)
  wire _05941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9815" *)
  wire _05942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9819" *)
  wire _05943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9820" *)
  wire _05944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9820" *)
  wire _05945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9820" *)
  wire _05946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9820" *)
  wire _05947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9823" *)
  wire _05948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9825" *)
  wire _05949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9825" *)
  wire _05950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9825" *)
  wire _05951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9830" *)
  wire _05952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9830" *)
  wire _05953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9832" *)
  wire _05954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9832" *)
  wire _05955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9833" *)
  wire _05956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9833" *)
  wire _05957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9837" *)
  wire _05958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9838" *)
  wire _05959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9838" *)
  wire _05960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9838" *)
  wire _05961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9838" *)
  wire _05962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9841" *)
  wire _05963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9843" *)
  wire _05964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9843" *)
  wire _05965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9843" *)
  wire _05966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9848" *)
  wire _05967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9848" *)
  wire _05968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9850" *)
  wire _05969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9850" *)
  wire _05970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9851" *)
  wire _05971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9851" *)
  wire _05972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9855" *)
  wire _05973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9856" *)
  wire _05974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9856" *)
  wire _05975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9856" *)
  wire _05976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9856" *)
  wire _05977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9859" *)
  wire _05978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9861" *)
  wire _05979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9861" *)
  wire _05980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9861" *)
  wire _05981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9866" *)
  wire _05982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9866" *)
  wire _05983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9868" *)
  wire _05984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9868" *)
  wire _05985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9869" *)
  wire _05986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9869" *)
  wire _05987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9873" *)
  wire _05988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9874" *)
  wire _05989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9874" *)
  wire _05990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9874" *)
  wire _05991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9874" *)
  wire _05992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9877" *)
  wire _05993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9879" *)
  wire _05994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9879" *)
  wire _05995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9879" *)
  wire _05996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9881" *)
  wire _05997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9886" *)
  wire _05998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9886" *)
  wire _05999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9886" *)
  wire _06000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9887" *)
  wire _06001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9890" *)
  wire _06002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9895" *)
  wire _06003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9895" *)
  wire _06004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9895" *)
  wire _06005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9896" *)
  wire _06006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9899" *)
  wire _06007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9904" *)
  wire _06008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9904" *)
  wire _06009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9904" *)
  wire _06010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9905" *)
  wire _06011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9910" *)
  wire _06012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9915" *)
  wire _06013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9915" *)
  wire _06014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9916" *)
  wire _06015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9916" *)
  wire _06016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *)
  wire _06017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *)
  wire _06018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *)
  wire _06019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *)
  wire _06020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *)
  wire _06021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *)
  wire _06022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *)
  wire _06023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *)
  wire _06024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *)
  wire [21:0] _06025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *)
  wire [21:0] _06026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *)
  wire [21:0] _06027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *)
  wire [21:0] _06028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *)
  wire [21:0] _06029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *)
  wire [21:0] _06030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *)
  wire [21:0] _06031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *)
  wire [21:0] _06032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *)
  wire [22:0] _06033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *)
  wire [22:0] _06034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *)
  wire [22:0] _06035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *)
  wire [22:0] _06036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *)
  wire [22:0] _06037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *)
  wire [22:0] _06038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *)
  wire [22:0] _06039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *)
  wire [22:0] _06040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *)
  wire [22:0] _06041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *)
  wire [22:0] _06042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *)
  wire [22:0] _06043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *)
  wire [22:0] _06044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *)
  wire [22:0] _06045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *)
  wire [22:0] _06046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *)
  wire [22:0] _06047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *)
  wire [22:0] _06048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *)
  wire [7:0] _06049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *)
  wire [7:0] _06050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *)
  wire [7:0] _06051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *)
  wire [7:0] _06052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3466" *)
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3462" *)
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3458" *)
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3454" *)
  wire FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3477" *)
  wire FpMantRNE_48U_24U_else_and_11_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3479" *)
  wire FpMantRNE_48U_24U_else_and_13_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3475" *)
  wire FpMantRNE_48U_24U_else_and_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3473" *)
  wire FpMantRNE_48U_24U_else_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2953" *)
  reg FpMantRNE_48U_24U_else_carry_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3022" *)
  reg FpMantRNE_48U_24U_else_carry_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3347" *)
  wire FpMantRNE_48U_24U_else_carry_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2959" *)
  reg FpMantRNE_48U_24U_else_carry_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3031" *)
  reg FpMantRNE_48U_24U_else_carry_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3354" *)
  wire FpMantRNE_48U_24U_else_carry_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2965" *)
  reg FpMantRNE_48U_24U_else_carry_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3040" *)
  reg FpMantRNE_48U_24U_else_carry_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3361" *)
  wire FpMantRNE_48U_24U_else_carry_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2971" *)
  reg FpMantRNE_48U_24U_else_carry_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3049" *)
  reg FpMantRNE_48U_24U_else_carry_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3368" *)
  wire FpMantRNE_48U_24U_else_carry_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4029" *)
  wire FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4033" *)
  wire FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4037" *)
  wire FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4041" *)
  wire FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3222" *)
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3218" *)
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3214" *)
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3210" *)
  wire FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3223" *)
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3219" *)
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3215" *)
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3211" *)
  wire [7:0] FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3993" *)
  wire [22:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4001" *)
  wire [22:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4009" *)
  wire [22:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4017" *)
  wire [22:0] FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3076" *)
  reg FpMul_8U_23U_FpMul_8U_23U_and_12_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3077" *)
  reg FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3355" *)
  wire FpMul_8U_23U_FpMul_8U_23U_and_12_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3095" *)
  reg FpMul_8U_23U_FpMul_8U_23U_and_13_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3096" *)
  reg FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3362" *)
  wire FpMul_8U_23U_FpMul_8U_23U_and_13_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3114" *)
  reg FpMul_8U_23U_FpMul_8U_23U_and_14_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3115" *)
  reg FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3369" *)
  wire FpMul_8U_23U_FpMul_8U_23U_and_14_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3522" *)
  wire [7:0] FpMul_8U_23U_FpMul_8U_23U_and_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3538" *)
  wire [7:0] FpMul_8U_23U_FpMul_8U_23U_and_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3554" *)
  wire [7:0] FpMul_8U_23U_FpMul_8U_23U_and_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3570" *)
  wire [7:0] FpMul_8U_23U_FpMul_8U_23U_and_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3057" *)
  reg FpMul_8U_23U_FpMul_8U_23U_and_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3058" *)
  reg FpMul_8U_23U_FpMul_8U_23U_and_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3348" *)
  wire FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4007" *)
  wire FpMul_8U_23U_FpMul_8U_23U_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4015" *)
  wire FpMul_8U_23U_FpMul_8U_23U_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4023" *)
  wire FpMul_8U_23U_FpMul_8U_23U_nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4027" *)
  wire FpMul_8U_23U_FpMul_8U_23U_nor_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3999" *)
  wire FpMul_8U_23U_FpMul_8U_23U_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4000" *)
  wire FpMul_8U_23U_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4008" *)
  wire FpMul_8U_23U_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4016" *)
  wire FpMul_8U_23U_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4024" *)
  wire FpMul_8U_23U_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3074" *)
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3075" *)
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3353" *)
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3093" *)
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3094" *)
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3360" *)
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3112" *)
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3113" *)
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3367" *)
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3055" *)
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3056" *)
  reg FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3346" *)
  wire FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3967" *)
  wire [7:0] FpMul_8U_23U_else_2_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3969" *)
  wire [7:0] FpMul_8U_23U_else_2_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3971" *)
  wire [7:0] FpMul_8U_23U_else_2_else_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3965" *)
  wire [7:0] FpMul_8U_23U_else_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3451" *)
  wire FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3054" *)
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3147" *)
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3073" *)
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3160" *)
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3092" *)
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3173" *)
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3111" *)
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3186" *)
  reg FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3208" *)
  wire FpMul_8U_23U_is_inf_1_lpi_1_dfm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3417" *)
  wire FpMul_8U_23U_lor_10_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3419" *)
  wire FpMul_8U_23U_lor_11_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3045" *)
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3046" *)
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3388" *)
  wire FpMul_8U_23U_lor_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3109" *)
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3181" *)
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3183" *)
  reg FpMul_8U_23U_lor_1_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3421" *)
  wire FpMul_8U_23U_lor_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3018" *)
  reg FpMul_8U_23U_lor_6_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3019" *)
  reg FpMul_8U_23U_lor_6_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3382" *)
  wire FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3052" *)
  reg FpMul_8U_23U_lor_6_lpi_1_dfm_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3142" *)
  reg FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3144" *)
  reg FpMul_8U_23U_lor_6_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3027" *)
  reg FpMul_8U_23U_lor_7_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3028" *)
  reg FpMul_8U_23U_lor_7_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3384" *)
  wire FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3071" *)
  reg FpMul_8U_23U_lor_7_lpi_1_dfm_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3155" *)
  reg FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3157" *)
  reg FpMul_8U_23U_lor_7_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3036" *)
  reg FpMul_8U_23U_lor_8_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3037" *)
  reg FpMul_8U_23U_lor_8_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3386" *)
  wire FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3090" *)
  reg FpMul_8U_23U_lor_8_lpi_1_dfm_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3168" *)
  reg FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3170" *)
  reg FpMul_8U_23U_lor_8_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3415" *)
  wire FpMul_8U_23U_lor_9_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3134" *)
  reg FpMul_8U_23U_mux_10_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3135" *)
  reg FpMul_8U_23U_mux_10_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3132" *)
  reg FpMul_8U_23U_mux_23_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3133" *)
  reg FpMul_8U_23U_mux_23_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3130" *)
  reg FpMul_8U_23U_mux_36_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3131" *)
  reg FpMul_8U_23U_mux_36_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3128" *)
  reg FpMul_8U_23U_mux_49_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3129" *)
  reg FpMul_8U_23U_mux_49_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4002" *)
  wire [22:0] FpMul_8U_23U_nor_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4010" *)
  wire [22:0] FpMul_8U_23U_nor_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4018" *)
  wire [22:0] FpMul_8U_23U_nor_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3994" *)
  wire [22:0] FpMul_8U_23U_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3221" *)
  wire [7:0] FpMul_8U_23U_o_expo_1_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3217" *)
  wire [7:0] FpMul_8U_23U_o_expo_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3213" *)
  wire [7:0] FpMul_8U_23U_o_expo_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3209" *)
  wire [7:0] FpMul_8U_23U_o_expo_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3398" *)
  wire [22:0] FpMul_8U_23U_o_mant_1_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3401" *)
  wire [22:0] FpMul_8U_23U_o_mant_2_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3404" *)
  wire [22:0] FpMul_8U_23U_o_mant_3_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3407" *)
  wire [22:0] FpMul_8U_23U_o_mant_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4048" *)
  wire [8:0] FpMul_8U_23U_oelse_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4052" *)
  wire [8:0] FpMul_8U_23U_oelse_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4056" *)
  wire [8:0] FpMul_8U_23U_oelse_1_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4044" *)
  wire [8:0] FpMul_8U_23U_oelse_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3484" *)
  wire FpMul_8U_23U_oelse_1_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3485" *)
  wire FpMul_8U_23U_oelse_1_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3486" *)
  wire FpMul_8U_23U_oelse_1_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3487" *)
  wire FpMul_8U_23U_oelse_1_and_7_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3892" *)
  wire FpMul_8U_23U_oelse_1_mux_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3903" *)
  wire FpMul_8U_23U_oelse_1_mux_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3914" *)
  wire FpMul_8U_23U_oelse_1_mux_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3925" *)
  wire FpMul_8U_23U_oelse_1_mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4028" *)
  wire FpMul_8U_23U_or_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4032" *)
  wire FpMul_8U_23U_or_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4036" *)
  wire FpMul_8U_23U_or_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4040" *)
  wire FpMul_8U_23U_or_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3414" *)
  wire [7:0] FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2952" *)
  reg [7:0] FpMul_8U_23U_p_expo_1_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3344" *)
  wire [7:0] FpMul_8U_23U_p_expo_1_sva_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3021" *)
  reg [7:0] FpMul_8U_23U_p_expo_1_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3416" *)
  wire [7:0] FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2958" *)
  reg [7:0] FpMul_8U_23U_p_expo_2_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3351" *)
  wire [7:0] FpMul_8U_23U_p_expo_2_sva_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3030" *)
  reg [7:0] FpMul_8U_23U_p_expo_2_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3418" *)
  wire [7:0] FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2964" *)
  reg [7:0] FpMul_8U_23U_p_expo_3_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3358" *)
  wire [7:0] FpMul_8U_23U_p_expo_3_sva_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3039" *)
  reg [7:0] FpMul_8U_23U_p_expo_3_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3461" *)
  wire FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3457" *)
  wire FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3453" *)
  wire FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3465" *)
  wire FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3285" *)
  wire FpMul_8U_23U_p_expo_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3288" *)
  wire FpMul_8U_23U_p_expo_and_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3292" *)
  wire FpMul_8U_23U_p_expo_and_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3281" *)
  wire FpMul_8U_23U_p_expo_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3420" *)
  wire [7:0] FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2970" *)
  reg [7:0] FpMul_8U_23U_p_expo_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3365" *)
  wire [7:0] FpMul_8U_23U_p_expo_sva_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3048" *)
  reg [7:0] FpMul_8U_23U_p_expo_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3314" *)
  wire [45:0] FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3315" *)
  wire [45:0] FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3316" *)
  wire [45:0] FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3317" *)
  wire [45:0] FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2951" *)
  reg [47:0] FpMul_8U_23U_p_mant_p1_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3232" *)
  wire [47:0] FpMul_8U_23U_p_mant_p1_1_sva_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2957" *)
  reg [47:0] FpMul_8U_23U_p_mant_p1_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3231" *)
  wire [47:0] FpMul_8U_23U_p_mant_p1_2_sva_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2963" *)
  reg [47:0] FpMul_8U_23U_p_mant_p1_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3230" *)
  wire [47:0] FpMul_8U_23U_p_mant_p1_3_sva_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3988" *)
  wire FpMul_8U_23U_p_mant_p1_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3983" *)
  wire FpMul_8U_23U_p_mant_p1_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3978" *)
  wire FpMul_8U_23U_p_mant_p1_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3973" *)
  wire FpMul_8U_23U_p_mant_p1_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2969" *)
  reg [47:0] FpMul_8U_23U_p_mant_p1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3229" *)
  wire [47:0] FpMul_8U_23U_p_mant_p1_sva_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3243" *)
  wire [64:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3202" *)
  reg [31:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3201" *)
  reg IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_64_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3241" *)
  wire [64:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3200" *)
  reg [31:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3199" *)
  reg IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_64_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3239" *)
  wire [64:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3198" *)
  reg [31:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3197" *)
  reg IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_64_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3237" *)
  wire [64:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3196" *)
  reg [31:0] IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3195" *)
  reg IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_64_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3449" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_10_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3450" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_11_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3474" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_13_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3476" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_16_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3478" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_19_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3480" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_22_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3287" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3290" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3294" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3447" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3448" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3283" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3400" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3403" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3406" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3409" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3228" *)
  wire [1086:0] IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3227" *)
  wire [1086:0] IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3226" *)
  wire [1086:0] IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3225" *)
  wire [1086:0] IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3399" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3402" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3405" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3408" *)
  wire IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3460" *)
  wire IsNaN_8U_23U_1_aelse_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3464" *)
  wire IsNaN_8U_23U_1_aelse_and_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3468" *)
  wire IsNaN_8U_23U_1_aelse_and_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3456" *)
  wire IsNaN_8U_23U_1_aelse_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3005" *)
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3006" *)
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3383" *)
  wire IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3000" *)
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3001" *)
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3385" *)
  wire IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2995" *)
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2996" *)
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3387" *)
  wire IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2990" *)
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2991" *)
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3389" *)
  wire IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2831" *)
  wire IsNaN_8U_23U_1_nor_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2830" *)
  wire IsNaN_8U_23U_1_nor_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2829" *)
  wire IsNaN_8U_23U_1_nor_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2832" *)
  wire IsNaN_8U_23U_1_nor_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3471" *)
  wire IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3455" *)
  wire IsNaN_8U_23U_aelse_and_17_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3459" *)
  wire IsNaN_8U_23U_aelse_and_19_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3463" *)
  wire IsNaN_8U_23U_aelse_and_21_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3467" *)
  wire IsNaN_8U_23U_aelse_and_23_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3470" *)
  wire IsNaN_8U_23U_aelse_and_24_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3481" *)
  wire IsNaN_8U_23U_aelse_and_25_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3482" *)
  wire IsNaN_8U_23U_aelse_and_26_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3483" *)
  wire IsNaN_8U_23U_aelse_and_27_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3296" *)
  wire IsNaN_8U_23U_aelse_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3297" *)
  wire IsNaN_8U_23U_aelse_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3298" *)
  wire IsNaN_8U_23U_aelse_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3299" *)
  wire IsNaN_8U_23U_aelse_and_7_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3279" *)
  wire IsNaN_8U_23U_aelse_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3002" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3003" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3004" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3394" *)
  wire IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3061" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3149" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3150" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3151" *)
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2997" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2998" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2999" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3395" *)
  wire IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3080" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3162" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3163" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3164" *)
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2992" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2993" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2994" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3396" *)
  wire IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3099" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3175" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3176" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3177" *)
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2987" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2988" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2989" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3397" *)
  wire IsNaN_8U_23U_land_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3118" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3188" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3189" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3190" *)
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2818" *)
  wire IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2817" *)
  wire IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2816" *)
  wire IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2819" *)
  wire IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3440" *)
  wire IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2949" *)
  reg IsZero_8U_23U_1_land_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3017" *)
  reg IsZero_8U_23U_1_land_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2955" *)
  reg IsZero_8U_23U_1_land_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3026" *)
  reg IsZero_8U_23U_1_land_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2961" *)
  reg IsZero_8U_23U_1_land_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3035" *)
  reg IsZero_8U_23U_1_land_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2967" *)
  reg IsZero_8U_23U_1_land_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3044" *)
  reg IsZero_8U_23U_1_land_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2948" *)
  reg IsZero_8U_23U_land_1_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3015" *)
  reg IsZero_8U_23U_land_1_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3016" *)
  reg IsZero_8U_23U_land_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3373" *)
  wire IsZero_8U_23U_land_1_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2954" *)
  reg IsZero_8U_23U_land_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3024" *)
  reg IsZero_8U_23U_land_2_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3025" *)
  reg IsZero_8U_23U_land_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3374" *)
  wire IsZero_8U_23U_land_2_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2960" *)
  reg IsZero_8U_23U_land_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3033" *)
  reg IsZero_8U_23U_land_3_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3034" *)
  reg IsZero_8U_23U_land_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3375" *)
  wire IsZero_8U_23U_land_3_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2966" *)
  reg IsZero_8U_23U_land_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3042" *)
  reg IsZero_8U_23U_land_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3043" *)
  reg IsZero_8U_23U_land_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3376" *)
  wire IsZero_8U_23U_land_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3446" *)
  wire MulIn_data_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3452" *)
  wire MulIn_data_and_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3280" *)
  wire MulIn_data_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3011" *)
  reg [127:0] MulIn_data_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3012" *)
  reg [127:0] MulIn_data_sva_132;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3013" *)
  reg [127:0] MulIn_data_sva_133;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3318" *)
  wire and_135_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3248" *)
  wire and_136_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3321" *)
  wire and_137_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3247" *)
  wire and_138_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3324" *)
  wire and_139_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3246" *)
  wire and_140_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3327" *)
  wire and_141_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3245" *)
  wire and_142_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3330" *)
  wire and_146_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3331" *)
  wire and_150_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3332" *)
  wire and_154_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3333" *)
  wire and_158_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2820" *)
  wire and_18_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2815" *)
  wire and_20_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3891" *)
  wire and_328_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3840" *)
  wire and_331_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3827" *)
  wire and_332_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3803" *)
  wire and_334_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3780" *)
  wire and_335_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3767" *)
  wire and_336_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3744" *)
  wire and_338_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3721" *)
  wire and_339_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3708" *)
  wire and_340_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3685" *)
  wire and_342_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3662" *)
  wire and_343_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3610" *)
  wire and_344_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3574" *)
  wire and_352_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3575" *)
  wire and_353_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3558" *)
  wire and_354_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3559" *)
  wire and_355_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3542" *)
  wire and_356_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3543" *)
  wire and_357_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3526" *)
  wire and_358_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3527" *)
  wire and_359_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3860" *)
  wire and_39_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3869" *)
  wire and_40_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3878" *)
  wire and_41_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2894" *)
  wire and_dcpl_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2895" *)
  wire and_dcpl_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2896" *)
  wire and_dcpl_24;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2897" *)
  wire and_dcpl_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2898" *)
  wire and_dcpl_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2886" *)
  wire and_dcpl_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2900" *)
  wire and_dcpl_30;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2902" *)
  wire and_dcpl_37;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2903" *)
  wire and_dcpl_38;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2904" *)
  wire and_dcpl_39;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2905" *)
  wire and_dcpl_45;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2906" *)
  wire and_dcpl_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2907" *)
  wire and_dcpl_47;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2908" *)
  wire and_dcpl_48;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2909" *)
  wire and_dcpl_50;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2910" *)
  wire and_dcpl_51;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2911" *)
  wire and_dcpl_52;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2912" *)
  wire and_dcpl_54;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2913" *)
  wire and_dcpl_55;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2914" *)
  wire and_dcpl_57;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2915" *)
  wire and_dcpl_58;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2888" *)
  wire and_dcpl_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2916" *)
  wire and_dcpl_60;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2917" *)
  wire and_dcpl_61;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2918" *)
  wire and_dcpl_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2919" *)
  wire and_dcpl_64;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2920" *)
  wire and_dcpl_66;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2921" *)
  wire and_dcpl_67;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2922" *)
  wire and_dcpl_69;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2923" *)
  wire and_dcpl_70;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2893" *)
  wire and_tmp_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3432" *)
  wire asn_156;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3433" *)
  wire asn_158;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3434" *)
  wire asn_160;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3435" *)
  wire asn_162;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3436" *)
  wire asn_164;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3437" *)
  wire asn_166;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3438" *)
  wire asn_168;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3439" *)
  wire asn_170;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2751" *)
  output cfg_mul_bypass_rsc_triosy_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2793" *)
  wire cfg_mul_bypass_rsc_triosy_obj_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2771" *)
  input cfg_mul_bypass_rsc_triosy_obj_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2776" *)
  output cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_pff;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2764" *)
  input cfg_mul_bypass_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3008" *)
  reg [31:0] cfg_mul_op_1_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2754" *)
  output cfg_mul_op_rsc_triosy_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2796" *)
  wire cfg_mul_op_rsc_triosy_obj_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2774" *)
  input cfg_mul_op_rsc_triosy_obj_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2767" *)
  input [31:0] cfg_mul_op_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2752" *)
  output cfg_mul_prelu_rsc_triosy_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2794" *)
  wire cfg_mul_prelu_rsc_triosy_obj_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2772" *)
  input cfg_mul_prelu_rsc_triosy_obj_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2765" *)
  input cfg_mul_prelu_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3007" *)
  reg cfg_mul_src_1_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3051" *)
  reg cfg_mul_src_1_sva_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3137" *)
  reg cfg_mul_src_1_sva_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3381" *)
  wire cfg_mul_src_1_sva_st_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2753" *)
  output cfg_mul_src_rsc_triosy_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2795" *)
  wire cfg_mul_src_rsc_triosy_obj_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2773" *)
  input cfg_mul_src_rsc_triosy_obj_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2766" *)
  input cfg_mul_src_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2756" *)
  input [1:0] cfg_precision;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3009" *)
  reg [9:0] cfg_truncate_1_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3010" *)
  reg [9:0] cfg_truncate_1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2755" *)
  output cfg_truncate_rsc_triosy_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2797" *)
  wire cfg_truncate_rsc_triosy_obj_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2775" *)
  input cfg_truncate_rsc_triosy_obj_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2768" *)
  input [9:0] cfg_truncate_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2747" *)
  output chn_mul_in_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2746" *)
  input chn_mul_in_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2745" *)
  input [127:0] chn_mul_in_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2780" *)
  wire chn_mul_in_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2783" *)
  wire [127:0] chn_mul_in_rsci_d_mxwt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2779" *)
  reg chn_mul_in_rsci_iswt0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2782" *)
  reg chn_mul_in_rsci_ld_core_psct;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3340" *)
  wire chn_mul_in_rsci_ld_core_psct_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2760" *)
  input chn_mul_in_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2761" *)
  output chn_mul_in_rsci_oswt_unreg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2781" *)
  wire chn_mul_in_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2750" *)
  output chn_mul_op_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2749" *)
  input chn_mul_op_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2748" *)
  input [127:0] chn_mul_op_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2786" *)
  wire chn_mul_op_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2789" *)
  wire [127:0] chn_mul_op_rsci_d_mxwt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2785" *)
  reg chn_mul_op_rsci_iswt0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2788" *)
  reg chn_mul_op_rsci_ld_core_psct;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3341" *)
  wire chn_mul_op_rsci_ld_core_psct_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2762" *)
  input chn_mul_op_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2763" *)
  output chn_mul_op_rsci_oswt_unreg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2787" *)
  wire chn_mul_op_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3253" *)
  wire chn_mul_out_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3254" *)
  wire chn_mul_out_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2759" *)
  output chn_mul_out_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2758" *)
  input chn_mul_out_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2757" *)
  output [127:0] chn_mul_out_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2791" *)
  wire chn_mul_out_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2813" *)
  reg chn_mul_out_rsci_d_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2800" *)
  reg [21:0] chn_mul_out_rsci_d_118_97;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2799" *)
  reg [7:0] chn_mul_out_rsci_d_126_119;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2798" *)
  reg chn_mul_out_rsci_d_127;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2812" *)
  reg [21:0] chn_mul_out_rsci_d_22_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2811" *)
  reg [7:0] chn_mul_out_rsci_d_30_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2810" *)
  reg chn_mul_out_rsci_d_31;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2809" *)
  reg chn_mul_out_rsci_d_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2808" *)
  reg [21:0] chn_mul_out_rsci_d_54_33;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2807" *)
  reg [7:0] chn_mul_out_rsci_d_62_55;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2806" *)
  reg chn_mul_out_rsci_d_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2805" *)
  reg chn_mul_out_rsci_d_64;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2804" *)
  reg [21:0] chn_mul_out_rsci_d_86_65;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2803" *)
  reg [7:0] chn_mul_out_rsci_d_94_87;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2802" *)
  reg chn_mul_out_rsci_d_95;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2801" *)
  reg chn_mul_out_rsci_d_96;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2790" *)
  reg chn_mul_out_rsci_iswt0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2769" *)
  input chn_mul_out_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2770" *)
  output chn_mul_out_rsci_oswt_unreg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2792" *)
  wire chn_mul_out_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2778" *)
  wire core_wen;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2784" *)
  wire core_wten;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3191" *)
  reg [30:0] else_MulOp_data_0_lpi_1_dfm_2_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3236" *)
  wire [30:0] else_MulOp_data_0_lpi_1_dfm_mx0_30_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3422" *)
  wire [31:0] else_MulOp_data_0_lpi_1_dfm_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3192" *)
  reg [30:0] else_MulOp_data_1_lpi_1_dfm_2_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3235" *)
  wire [30:0] else_MulOp_data_1_lpi_1_dfm_mx0_30_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3423" *)
  wire [31:0] else_MulOp_data_1_lpi_1_dfm_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3193" *)
  reg [30:0] else_MulOp_data_2_lpi_1_dfm_2_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3234" *)
  wire [30:0] else_MulOp_data_2_lpi_1_dfm_mx0_30_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3424" *)
  wire [31:0] else_MulOp_data_2_lpi_1_dfm_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3194" *)
  reg [30:0] else_MulOp_data_3_lpi_1_dfm_2_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3233" *)
  wire [30:0] else_MulOp_data_3_lpi_1_dfm_mx0_30_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3425" *)
  wire [31:0] else_MulOp_data_3_lpi_1_dfm_mx1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3443" *)
  wire else_MulOp_data_and_10_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3444" *)
  wire else_MulOp_data_and_11_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3282" *)
  wire else_MulOp_data_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3286" *)
  wire else_MulOp_data_and_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3289" *)
  wire else_MulOp_data_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3293" *)
  wire else_MulOp_data_and_7_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3441" *)
  wire else_MulOp_data_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3442" *)
  wire else_MulOp_data_and_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3063" *)
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3064" *)
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3062" *)
  reg [7:0] else_MulOp_data_slc_else_MulOp_data_0_30_23_5_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3082" *)
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3083" *)
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3081" *)
  reg [7:0] else_MulOp_data_slc_else_MulOp_data_1_30_23_5_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3101" *)
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3102" *)
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3100" *)
  reg [7:0] else_MulOp_data_slc_else_MulOp_data_2_30_23_5_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3120" *)
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3121" *)
  reg [22:0] else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3119" *)
  reg [7:0] else_MulOp_data_slc_else_MulOp_data_3_30_23_5_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3205" *)
  wire [7:0] else_mux_1_tmp_30_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3204" *)
  wire [7:0] else_mux_2_tmp_30_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3203" *)
  wire [7:0] else_mux_3_tmp_30_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3206" *)
  wire [7:0] else_mux_tmp_30_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2814" *)
  wire [1:0] fsm_output;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3014" *)
  reg io_read_cfg_mul_bypass_rsc_svs_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3136" *)
  reg io_read_cfg_mul_bypass_rsc_svs_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3139" *)
  reg io_read_cfg_mul_bypass_rsc_svs_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2972" *)
  reg main_stage_v_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3372" *)
  wire main_stage_v_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2973" *)
  reg main_stage_v_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3342" *)
  wire main_stage_v_2_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2974" *)
  reg main_stage_v_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3343" *)
  wire main_stage_v_3_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3996" *)
  wire [22:0] mul_mul_1_FpMantRNE_48U_24U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3023" *)
  reg mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3060" *)
  reg mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3148" *)
  reg mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2828" *)
  wire mul_mul_1_FpMantRNE_48U_24U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3059" *)
  reg [22:0] mul_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3976" *)
  (* unused_bits = "0" *)
  wire [8:0] mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3496" *)
  wire mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4062" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4025" *)
  wire [7:0] mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3053" *)
  reg mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3146" *)
  reg mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3488" *)
  wire mul_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3974" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2950" *)
  reg mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3020" *)
  reg mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3143" *)
  reg mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3145" *)
  reg mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3492" *)
  wire mul_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4042" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8" *)
  wire [9:0] mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2824" *)
  wire [47:0] mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3899" *)
  wire mul_mul_1_FpMul_8U_23U_xor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3065" *)
  reg [63:0] mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3066" *)
  reg [63:0] mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3390" *)
  wire [63:0] mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3518" *)
  wire mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3531" *)
  wire mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3524" *)
  wire [7:0] mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3519" *)
  wire [21:0] mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4058" *)
  wire mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3069" *)
  reg mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3070" *)
  reg mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3349" *)
  wire mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3067" *)
  reg mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3068" *)
  reg mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3350" *)
  wire mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3520" *)
  wire [21:0] mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3525" *)
  wire [7:0] mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4004" *)
  wire [22:0] mul_mul_2_FpMantRNE_48U_24U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3032" *)
  reg mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3079" *)
  reg mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3161" *)
  reg mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2827" *)
  wire mul_mul_2_FpMantRNE_48U_24U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3078" *)
  reg [22:0] mul_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3981" *)
  (* unused_bits = "0" *)
  wire [8:0] mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3497" *)
  wire mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4066" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4030" *)
  wire [7:0] mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3072" *)
  reg mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3159" *)
  reg mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3489" *)
  wire mul_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3979" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2956" *)
  reg mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3029" *)
  reg mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3156" *)
  reg mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3158" *)
  reg mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3493" *)
  wire mul_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4046" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8" *)
  wire [9:0] mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2823" *)
  wire [47:0] mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3910" *)
  wire mul_mul_2_FpMul_8U_23U_xor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3084" *)
  reg [63:0] mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3085" *)
  reg [63:0] mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3391" *)
  wire [63:0] mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3534" *)
  wire mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3547" *)
  wire mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3540" *)
  wire [7:0] mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3535" *)
  wire [21:0] mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4059" *)
  wire mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3088" *)
  reg mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3089" *)
  reg mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3356" *)
  wire mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3086" *)
  reg mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3087" *)
  reg mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3357" *)
  wire mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3536" *)
  wire [21:0] mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3541" *)
  wire [7:0] mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4012" *)
  wire [22:0] mul_mul_3_FpMantRNE_48U_24U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3041" *)
  reg mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3098" *)
  reg mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3174" *)
  reg mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2826" *)
  wire mul_mul_3_FpMantRNE_48U_24U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3097" *)
  reg [22:0] mul_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3986" *)
  (* unused_bits = "0" *)
  wire [8:0] mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3498" *)
  wire mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4070" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4034" *)
  wire [7:0] mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3091" *)
  reg mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3172" *)
  reg mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3490" *)
  wire mul_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3984" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2962" *)
  reg mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3038" *)
  reg mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3169" *)
  reg mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3171" *)
  reg mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3494" *)
  wire mul_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4050" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8" *)
  wire [9:0] mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2822" *)
  wire [47:0] mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3921" *)
  wire mul_mul_3_FpMul_8U_23U_xor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3103" *)
  reg [63:0] mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3104" *)
  reg [63:0] mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3392" *)
  wire [63:0] mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3550" *)
  wire mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3563" *)
  wire mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3556" *)
  wire [7:0] mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3551" *)
  wire [21:0] mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4060" *)
  wire mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3107" *)
  reg mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3108" *)
  reg mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3363" *)
  wire mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3105" *)
  reg mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3106" *)
  reg mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3364" *)
  wire mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3552" *)
  wire [21:0] mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3557" *)
  wire [7:0] mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4020" *)
  wire [22:0] mul_mul_4_FpMantRNE_48U_24U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3050" *)
  reg mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3117" *)
  reg mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3187" *)
  reg mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2825" *)
  wire mul_mul_4_FpMantRNE_48U_24U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3116" *)
  reg [22:0] mul_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3991" *)
  (* unused_bits = "0" *)
  wire [8:0] mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3499" *)
  wire mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4074" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4038" *)
  wire [7:0] mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3110" *)
  reg mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3185" *)
  reg mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3491" *)
  wire mul_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3989" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2968" *)
  reg mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3047" *)
  reg mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3182" *)
  reg mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3184" *)
  reg mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3495" *)
  wire mul_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4054" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8" *)
  wire [9:0] mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2821" *)
  wire [47:0] mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3932" *)
  wire mul_mul_4_FpMul_8U_23U_xor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3122" *)
  reg [63:0] mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3123" *)
  reg [63:0] mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3393" *)
  wire [63:0] mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3566" *)
  wire mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3579" *)
  wire mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3572" *)
  wire [7:0] mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3567" *)
  wire [21:0] mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4061" *)
  wire mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3126" *)
  reg mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3127" *)
  reg mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3370" *)
  wire mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3124" *)
  reg mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3125" *)
  reg mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3371" *)
  wire mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3568" *)
  wire [21:0] mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3573" *)
  wire [7:0] mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3469" *)
  wire mul_mul_aelse_and_12_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3472" *)
  wire mul_mul_aelse_and_19_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3445" *)
  wire mul_mul_aelse_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3251" *)
  wire mul_mul_and_17_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3250" *)
  wire mul_mul_and_19_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3249" *)
  wire mul_mul_and_21_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3252" *)
  wire mul_mul_and_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3578" *)
  wire mul_mul_else_mux_104_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3565" *)
  wire mul_mul_else_mux_107_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3530" *)
  wire mul_mul_else_mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3517" *)
  wire mul_mul_else_mux_26_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3546" *)
  wire mul_mul_else_mux_50_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3533" *)
  wire mul_mul_else_mux_53_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3562" *)
  wire mul_mul_else_mux_77_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3549" *)
  wire mul_mul_else_mux_80_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3207" *)
  wire mul_mul_else_unequal_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3329" *)
  wire mul_mul_if_and_1_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3325" *)
  wire mul_mul_if_and_2_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3326" *)
  wire mul_mul_if_and_3_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3322" *)
  wire mul_mul_if_and_4_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3323" *)
  wire mul_mul_if_and_5_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3319" *)
  wire mul_mul_if_and_6_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3320" *)
  wire mul_mul_if_and_7_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3328" *)
  wire mul_mul_if_and_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2975" *)
  reg mul_mul_land_1_lpi_1_dfm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2976" *)
  reg mul_mul_land_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2977" *)
  reg mul_mul_land_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3380" *)
  wire mul_mul_land_1_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3138" *)
  reg mul_mul_land_1_lpi_1_dfm_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3140" *)
  reg mul_mul_land_1_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3141" *)
  reg mul_mul_land_1_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2978" *)
  reg mul_mul_land_2_lpi_1_dfm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2979" *)
  reg mul_mul_land_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2980" *)
  reg mul_mul_land_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3379" *)
  wire mul_mul_land_2_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3152" *)
  reg mul_mul_land_2_lpi_1_dfm_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3153" *)
  reg mul_mul_land_2_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3154" *)
  reg mul_mul_land_2_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2981" *)
  reg mul_mul_land_3_lpi_1_dfm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2982" *)
  reg mul_mul_land_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2983" *)
  reg mul_mul_land_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3378" *)
  wire mul_mul_land_3_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3165" *)
  reg mul_mul_land_3_lpi_1_dfm_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3166" *)
  reg mul_mul_land_3_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3167" *)
  reg mul_mul_land_3_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2984" *)
  reg mul_mul_land_lpi_1_dfm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2985" *)
  reg mul_mul_land_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2986" *)
  reg mul_mul_land_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3377" *)
  wire mul_mul_land_lpi_1_dfm_mx1w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3178" *)
  reg mul_mul_land_lpi_1_dfm_st_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3179" *)
  reg mul_mul_land_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3180" *)
  reg mul_mul_land_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3412" *)
  wire mul_mul_mul_mul_nor_2_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3411" *)
  wire mul_mul_mul_mul_nor_4_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3410" *)
  wire mul_mul_mul_mul_nor_6_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3413" *)
  wire mul_mul_mul_mul_nor_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3516" *)
  wire mul_mul_mux_108_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3529" *)
  wire mul_mul_mux_109_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3532" *)
  wire mul_mul_mux_110_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3545" *)
  wire mul_mul_mux_111_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3548" *)
  wire mul_mul_mux_112_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3561" *)
  wire mul_mul_mux_113_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3564" *)
  wire mul_mul_mux_114_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3577" *)
  wire mul_mul_mux_115_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3737" *)
  wire mux_100_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3731" *)
  wire mux_101_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3729" *)
  wire mux_102_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3742" *)
  wire mux_103_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3740" *)
  wire mux_104_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3727" *)
  wire mux_105_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3746" *)
  wire mux_106_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3745" *)
  wire mux_107_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3754" *)
  wire mux_108_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3753" *)
  wire mux_109_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4083" *)
  wire mux_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3757" *)
  wire mux_110_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3752" *)
  wire mux_111_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3750" *)
  wire mux_112_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3760" *)
  wire mux_113_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3765" *)
  wire mux_115_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3763" *)
  wire mux_116_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4119" *)
  wire mux_117_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4117" *)
  wire mux_118_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3773" *)
  wire mux_121_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3771" *)
  wire mux_122_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3768" *)
  wire mux_123_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3766" *)
  wire mux_124_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3339" *)
  wire mux_125_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3781" *)
  wire mux_126_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3779" *)
  wire mux_127_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3778" *)
  wire mux_128_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3792" *)
  wire mux_129_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3335" *)
  wire mux_12_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3791" *)
  wire mux_130_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3796" *)
  wire mux_131_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3790" *)
  wire mux_132_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3788" *)
  wire mux_133_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3801" *)
  wire mux_134_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3799" *)
  wire mux_135_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3786" *)
  wire mux_136_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3805" *)
  wire mux_137_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3804" *)
  wire mux_138_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3813" *)
  wire mux_139_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3585" *)
  wire mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3812" *)
  wire mux_140_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3816" *)
  wire mux_141_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3811" *)
  wire mux_142_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3809" *)
  wire mux_143_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4124" *)
  wire mux_144_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3821" *)
  wire mux_146_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3819" *)
  wire mux_147_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3825" *)
  wire mux_148_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3823" *)
  wire mux_149_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3584" *)
  wire mux_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4127" *)
  wire mux_150_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3833" *)
  wire mux_153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3831" *)
  wire mux_154_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3828" *)
  wire mux_155_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3826" *)
  wire mux_156_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3841" *)
  wire mux_157_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3839" *)
  wire mux_158_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3838" *)
  wire mux_159_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4088" *)
  wire mux_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3846" *)
  wire mux_160_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3939" *)
  wire mux_161_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3938" *)
  wire mux_162_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3937" *)
  wire mux_163_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3936" *)
  wire mux_164_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3848" *)
  wire mux_168_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3946" *)
  wire mux_169_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3945" *)
  wire mux_170_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3944" *)
  wire mux_171_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3943" *)
  wire mux_172_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3850" *)
  wire mux_173_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3953" *)
  wire mux_174_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3952" *)
  wire mux_175_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3951" *)
  wire mux_176_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3950" *)
  wire mux_177_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3852" *)
  wire mux_178_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3961" *)
  wire mux_179_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3336" *)
  wire mux_17_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3960" *)
  wire mux_180_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3959" *)
  wire mux_181_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3957" *)
  wire mux_182_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3855" *)
  wire mux_184_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3854" *)
  wire mux_185_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3861" *)
  wire mux_186_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3859" *)
  wire mux_187_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3865" *)
  wire mux_188_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3864" *)
  wire mux_189_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3589" *)
  wire mux_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3870" *)
  wire mux_190_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3868" *)
  wire mux_191_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3874" *)
  wire mux_192_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3873" *)
  wire mux_193_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3879" *)
  wire mux_194_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3877" *)
  wire mux_195_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3883" *)
  wire mux_196_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3882" *)
  wire mux_197_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3888" *)
  wire mux_198_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3890" *)
  wire mux_199_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3588" *)
  wire mux_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3887" *)
  wire mux_200_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3886" *)
  wire mux_201_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3894" *)
  wire mux_202_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3893" *)
  wire mux_203_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3900" *)
  wire mux_207_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3905" *)
  wire mux_208_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3904" *)
  wire mux_209_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4092" *)
  wire mux_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3911" *)
  wire mux_213_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3916" *)
  wire mux_214_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3915" *)
  wire mux_215_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3922" *)
  wire mux_219_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3927" *)
  wire mux_220_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3926" *)
  wire mux_221_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3933" *)
  wire mux_225_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3337" *)
  wire mux_22_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4064" *)
  wire mux_233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4068" *)
  wire mux_234_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4072" *)
  wire mux_235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4076" *)
  wire mux_236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3995" *)
  wire [22:0] mux_237_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4003" *)
  wire [22:0] mux_238_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4011" *)
  wire [22:0] mux_239_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3593" *)
  wire mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4019" *)
  wire [22:0] mux_240_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3592" *)
  wire mux_24_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3596" *)
  wire mux_26_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3597" *)
  wire mux_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3600" *)
  wire mux_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3603" *)
  wire mux_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3606" *)
  wire mux_33_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3616" *)
  wire mux_35_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3615" *)
  wire mux_36_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3620" *)
  wire mux_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3614" *)
  wire mux_38_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3611" *)
  wire mux_39_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3625" *)
  wire mux_40_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3623" *)
  wire mux_41_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3609" *)
  wire mux_42_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3628" *)
  wire mux_43_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3627" *)
  wire mux_44_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3636" *)
  wire mux_45_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3635" *)
  wire mux_46_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3639" *)
  wire mux_47_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3634" *)
  wire mux_48_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3632" *)
  wire mux_49_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3642" *)
  wire mux_50_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4098" *)
  wire mux_52_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3647" *)
  wire mux_54_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3645" *)
  wire mux_55_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4102" *)
  wire mux_56_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4100" *)
  wire mux_57_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4078" *)
  wire mux_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3655" *)
  wire mux_60_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3653" *)
  wire mux_61_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3651" *)
  wire mux_62_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3649" *)
  wire mux_63_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3663" *)
  wire mux_64_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3661" *)
  wire mux_65_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3660" *)
  wire mux_66_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3674" *)
  wire mux_67_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3673" *)
  wire mux_68_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3678" *)
  wire mux_69_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3672" *)
  wire mux_70_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3670" *)
  wire mux_71_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3683" *)
  wire mux_72_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3681" *)
  wire mux_73_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3668" *)
  wire mux_74_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3687" *)
  wire mux_75_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3686" *)
  wire mux_76_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3695" *)
  wire mux_77_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3694" *)
  wire mux_78_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3698" *)
  wire mux_79_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3334" *)
  wire mux_7_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3693" *)
  wire mux_80_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3691" *)
  wire mux_81_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3701" *)
  wire mux_82_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3706" *)
  wire mux_84_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3704" *)
  wire mux_85_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4111" *)
  wire mux_86_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4109" *)
  wire mux_87_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3581" *)
  wire mux_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3714" *)
  wire mux_90_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3712" *)
  wire mux_91_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3709" *)
  wire mux_92_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3707" *)
  wire mux_93_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3338" *)
  wire mux_94_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3722" *)
  wire mux_95_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3720" *)
  wire mux_96_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3719" *)
  wire mux_97_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3733" *)
  wire mux_98_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3732" *)
  wire mux_99_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3580" *)
  wire mux_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2873" *)
  wire mux_tmp_109;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2882" *)
  wire mux_tmp_140;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2856" *)
  wire mux_tmp_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2857" *)
  wire mux_tmp_48;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2865" *)
  wire mux_tmp_78;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3654" *)
  wire nand_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3682" *)
  wire nand_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3713" *)
  wire nand_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3741" *)
  wire nand_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3772" *)
  wire nand_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3800" *)
  wire nand_34_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3832" *)
  wire nand_36_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3305" *)
  wire nand_42_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3304" *)
  wire nand_45_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3303" *)
  wire nand_48_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3224" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3220" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3216" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3212" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3968" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMul_8U_23U_else_2_else_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3970" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMul_8U_23U_else_2_else_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3972" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMul_8U_23U_else_2_else_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3966" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMul_8U_23U_else_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4049" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_FpMul_8U_23U_oelse_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4053" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_FpMul_8U_23U_oelse_1_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4057" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_FpMul_8U_23U_oelse_1_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4045" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_FpMul_8U_23U_oelse_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3345" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMul_8U_23U_p_expo_1_sva_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3352" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMul_8U_23U_p_expo_2_sva_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3359" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMul_8U_23U_p_expo_3_sva_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3366" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpMul_8U_23U_p_expo_sva_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3244" *)
  (* unused_bits = "65" *)
  wire [65:0] nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3242" *)
  (* unused_bits = "65" *)
  wire [65:0] nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3240" *)
  (* unused_bits = "65" *)
  wire [65:0] nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3238" *)
  (* unused_bits = "65" *)
  wire [65:0] nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4153" *)
  wire [127:0] nl_Y_mul_core_chn_mul_out_rsci_inst_chn_mul_out_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3997" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_mul_mul_1_FpMantRNE_48U_24U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3977" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4063" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4026" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3975" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4043" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 10" *)
  wire [10:0] nl_mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4133" *)
  wire [1086:0] nl_mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4136" *)
  wire [9:0] nl_mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4005" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_mul_mul_2_FpMantRNE_48U_24U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3982" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4067" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4031" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3980" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4047" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 10" *)
  wire [10:0] nl_mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4138" *)
  wire [1086:0] nl_mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4141" *)
  wire [9:0] nl_mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4013" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_mul_mul_3_FpMantRNE_48U_24U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3987" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4071" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4035" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3985" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4051" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 10" *)
  wire [10:0] nl_mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4143" *)
  wire [1086:0] nl_mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4146" *)
  wire [9:0] nl_mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4021" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_mul_mul_4_FpMantRNE_48U_24U_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3992" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4075" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4039" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3990" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9" *)
  wire [9:0] nl_mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4055" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 10" *)
  wire [10:0] nl_mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4148" *)
  wire [1086:0] nl_mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4151" *)
  wire [9:0] nl_mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3309" *)
  wire nor_115_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3308" *)
  wire nor_116_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3307" *)
  wire nor_117_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3306" *)
  wire nor_118_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3934" *)
  wire nor_119_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3935" *)
  wire nor_120_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3928" *)
  wire nor_121_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3929" *)
  wire nor_122_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3931" *)
  wire nor_123_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3923" *)
  wire nor_124_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3924" *)
  wire nor_125_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3917" *)
  wire nor_126_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3918" *)
  wire nor_127_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3920" *)
  wire nor_128_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3912" *)
  wire nor_129_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3913" *)
  wire nor_130_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3906" *)
  wire nor_131_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3907" *)
  wire nor_132_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3909" *)
  wire nor_133_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3901" *)
  wire nor_134_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3902" *)
  wire nor_135_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3895" *)
  wire nor_136_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3896" *)
  wire nor_137_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3898" *)
  wire nor_138_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3876" *)
  wire nor_140_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3867" *)
  wire nor_142_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3284" *)
  wire nor_143_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3857" *)
  wire nor_144_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3962" *)
  wire nor_153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3954" *)
  wire nor_155_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3947" *)
  wire nor_157_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3940" *)
  wire nor_159_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3842" *)
  wire nor_161_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3843" *)
  wire nor_163_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3844" *)
  wire nor_164_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3845" *)
  wire nor_165_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3829" *)
  wire nor_167_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3830" *)
  wire nor_168_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3834" *)
  wire nor_169_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3275" *)
  wire nor_170_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3835" *)
  wire nor_171_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3837" *)
  wire nor_172_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3277" *)
  wire nor_174_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4130" *)
  wire nor_175_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4131" *)
  wire nor_176_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4126" *)
  wire nor_177_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4128" *)
  wire nor_179_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4129" *)
  wire nor_180_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3810" *)
  wire nor_181_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3818" *)
  wire nor_183_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3806" *)
  wire nor_186_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3807" *)
  wire nor_187_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3808" *)
  wire nor_188_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3787" *)
  wire nor_189_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3273" *)
  wire nor_190_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3798" *)
  wire nor_192_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3274" *)
  wire nor_193_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3802" *)
  wire nor_194_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3782" *)
  wire nor_195_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3783" *)
  wire nor_197_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3784" *)
  wire nor_198_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3785" *)
  wire nor_199_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3553" *)
  wire nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3769" *)
  wire nor_201_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3770" *)
  wire nor_202_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3774" *)
  wire nor_203_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3270" *)
  wire nor_204_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3775" *)
  wire nor_205_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3777" *)
  wire nor_206_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3272" *)
  wire nor_208_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4122" *)
  wire nor_209_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4123" *)
  wire nor_210_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4116" *)
  wire nor_211_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4118" *)
  wire nor_212_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4120" *)
  wire nor_214_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4121" *)
  wire nor_215_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3761" *)
  wire nor_216_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3762" *)
  wire nor_217_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3751" *)
  wire nor_218_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3759" *)
  wire nor_220_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3747" *)
  wire nor_223_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3748" *)
  wire nor_224_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3749" *)
  wire nor_225_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3728" *)
  wire nor_226_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3268" *)
  wire nor_227_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3739" *)
  wire nor_229_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3269" *)
  wire nor_230_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3743" *)
  wire nor_231_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3723" *)
  wire nor_232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3724" *)
  wire nor_234_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3725" *)
  wire nor_235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3726" *)
  wire nor_236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3710" *)
  wire nor_238_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3711" *)
  wire nor_239_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3715" *)
  wire nor_240_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3265" *)
  wire nor_241_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3716" *)
  wire nor_242_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3718" *)
  wire nor_243_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3267" *)
  wire nor_245_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4114" *)
  wire nor_246_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4115" *)
  wire nor_247_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4108" *)
  wire nor_248_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4110" *)
  wire nor_249_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4112" *)
  wire nor_251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4113" *)
  wire nor_252_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3702" *)
  wire nor_253_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3703" *)
  wire nor_254_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3692" *)
  wire nor_255_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3700" *)
  wire nor_257_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3688" *)
  wire nor_260_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3689" *)
  wire nor_261_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3690" *)
  wire nor_262_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3669" *)
  wire nor_263_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3263" *)
  wire nor_264_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3680" *)
  wire nor_266_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3264" *)
  wire nor_267_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3684" *)
  wire nor_268_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3664" *)
  wire nor_269_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3665" *)
  wire nor_271_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3666" *)
  wire nor_272_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3667" *)
  wire nor_273_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3650" *)
  wire nor_275_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3656" *)
  wire nor_276_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3260" *)
  wire nor_277_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3657" *)
  wire nor_278_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3659" *)
  wire nor_279_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3262" *)
  wire nor_282_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4106" *)
  wire nor_283_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4107" *)
  wire nor_284_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4099" *)
  wire nor_285_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4101" *)
  wire nor_286_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4103" *)
  wire nor_288_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4104" *)
  wire nor_289_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3643" *)
  wire nor_290_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3644" *)
  wire nor_291_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3633" *)
  wire nor_292_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3641" *)
  wire nor_294_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3629" *)
  wire nor_296_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3630" *)
  wire nor_297_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3631" *)
  wire nor_298_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3612" *)
  wire nor_299_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3537" *)
  wire nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3613" *)
  wire nor_300_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3259" *)
  wire nor_301_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3622" *)
  wire nor_303_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3626" *)
  wire nor_304_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3607" *)
  wire nor_307_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3608" *)
  wire nor_308_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3604" *)
  wire nor_311_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3605" *)
  wire nor_312_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3601" *)
  wire nor_315_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3602" *)
  wire nor_316_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3598" *)
  wire nor_319_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3599" *)
  wire nor_320_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4093" *)
  wire nor_321_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4094" *)
  wire nor_322_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4095" *)
  wire nor_323_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4087" *)
  wire nor_324_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4090" *)
  wire nor_325_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4082" *)
  wire nor_326_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4085" *)
  wire nor_327_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4080" *)
  wire nor_331_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3885" *)
  wire nor_342_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3313" *)
  wire nor_346_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3312" *)
  wire nor_347_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3311" *)
  wire nor_348_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3521" *)
  wire nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3569" *)
  wire nor_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4077" *)
  wire nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2874" *)
  wire not_tmp_106;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2875" *)
  wire not_tmp_107;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2840" *)
  wire not_tmp_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2878" *)
  wire not_tmp_121;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2883" *)
  wire not_tmp_129;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2884" *)
  wire not_tmp_130;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2842" *)
  wire not_tmp_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2834" *)
  wire not_tmp_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2858" *)
  wire not_tmp_54;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2859" *)
  wire not_tmp_55;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2837" *)
  wire not_tmp_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2866" *)
  wire not_tmp_81;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2867" *)
  wire not_tmp_82;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2743" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2744" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3426" *)
  wire or_11_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3427" *)
  wire or_12_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3428" *)
  wire or_13_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3617" *)
  wire or_142_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3618" *)
  wire or_143_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3621" *)
  wire or_147_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3429" *)
  wire or_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3624" *)
  wire or_153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3430" *)
  wire or_15_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3637" *)
  wire or_165_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3638" *)
  wire or_166_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3640" *)
  wire or_169_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3431" *)
  wire or_16_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3646" *)
  wire or_181_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3648" *)
  wire or_185_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4097" *)
  wire or_187_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3310" *)
  wire or_189_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4105" *)
  wire or_193_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4079" *)
  wire or_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3658" *)
  wire or_210_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3652" *)
  wire or_211_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3671" *)
  wire or_227_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3675" *)
  wire or_230_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3676" *)
  wire or_231_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3679" *)
  wire or_235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3696" *)
  wire or_254_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3697" *)
  wire or_255_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3699" *)
  wire or_258_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4081" *)
  wire or_26_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3705" *)
  wire or_270_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3256" *)
  wire or_27_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3582" *)
  wire or_28_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3717" *)
  wire or_292_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3730" *)
  wire or_307_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3734" *)
  wire or_310_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3735" *)
  wire or_311_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3738" *)
  wire or_315_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3583" *)
  wire or_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3755" *)
  wire or_334_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3756" *)
  wire or_335_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3758" *)
  wire or_338_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4084" *)
  wire or_34_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3764" *)
  wire or_350_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3776" *)
  wire or_372_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3789" *)
  wire or_387_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3793" *)
  wire or_390_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3794" *)
  wire or_391_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3797" *)
  wire or_395_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4086" *)
  wire or_40_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3814" *)
  wire or_414_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3815" *)
  wire or_415_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3817" *)
  wire or_418_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3822" *)
  wire or_424_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3820" *)
  wire or_429_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3586" *)
  wire or_42_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3291" *)
  wire or_430_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4125" *)
  wire or_435_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3824" *)
  wire or_436_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3836" *)
  wire or_453_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3587" *)
  wire or_45_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3847" *)
  wire or_467_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3295" *)
  wire or_468_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3300" *)
  wire or_469_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3941" *)
  wire or_473_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3942" *)
  wire or_474_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3849" *)
  wire or_480_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3301" *)
  wire or_482_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3948" *)
  wire or_486_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3949" *)
  wire or_487_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3851" *)
  wire or_488_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4089" *)
  wire or_48_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3302" *)
  wire or_490_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3955" *)
  wire or_494_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3956" *)
  wire or_495_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3853" *)
  wire or_496_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3958" *)
  wire or_498_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3963" *)
  wire or_502_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3964" *)
  wire or_503_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3858" *)
  wire or_509_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3856" *)
  wire or_511_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3862" *)
  wire or_515_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3866" *)
  wire or_519_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3871" *)
  wire or_523_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3875" *)
  wire or_527_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3880" *)
  wire or_531_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3884" *)
  wire or_535_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3897" *)
  wire or_540_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4091" *)
  wire or_54_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3908" *)
  wire or_551_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3919" *)
  wire or_561_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3590" *)
  wire or_56_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3930" *)
  wire or_571_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3591" *)
  wire or_59_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4096" *)
  wire or_65_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3594" *)
  wire or_67_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3595" *)
  wire or_70_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4065" *)
  wire or_743_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4069" *)
  wire or_744_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4073" *)
  wire or_745_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3257" *)
  wire or_74_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3795" *)
  wire or_828_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3736" *)
  wire or_829_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3677" *)
  wire or_830_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3619" *)
  wire or_831_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3576" *)
  wire or_836_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3560" *)
  wire or_837_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3544" *)
  wire or_838_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3528" *)
  wire or_839_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4006" *)
  wire or_840_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4014" *)
  wire or_841_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4022" *)
  wire or_842_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2940" *)
  wire or_dcpl_102;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2941" *)
  wire or_dcpl_105;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2942" *)
  wire or_dcpl_108;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2943" *)
  wire or_dcpl_110;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2944" *)
  wire or_dcpl_125;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2901" *)
  wire or_dcpl_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2924" *)
  wire or_dcpl_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2925" *)
  wire or_dcpl_23;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2926" *)
  wire or_dcpl_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2927" *)
  wire or_dcpl_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2928" *)
  wire or_dcpl_37;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2929" *)
  wire or_dcpl_40;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2930" *)
  wire or_dcpl_50;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2931" *)
  wire or_dcpl_53;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2932" *)
  wire or_dcpl_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2933" *)
  wire or_dcpl_66;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2934" *)
  wire or_dcpl_75;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2899" *)
  wire or_dcpl_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2935" *)
  wire or_dcpl_81;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2936" *)
  wire or_dcpl_87;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2937" *)
  wire or_dcpl_93;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2938" *)
  wire or_dcpl_96;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2939" *)
  wire or_dcpl_99;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3998" *)
  wire or_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2833" *)
  wire or_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2848" *)
  wire or_tmp_107;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2835" *)
  wire or_tmp_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2849" *)
  wire or_tmp_123;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2850" *)
  wire or_tmp_128;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2851" *)
  wire or_tmp_132;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2852" *)
  wire or_tmp_133;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2853" *)
  wire or_tmp_146;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2836" *)
  wire or_tmp_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2854" *)
  wire or_tmp_167;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2855" *)
  wire or_tmp_173;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2860" *)
  wire or_tmp_211;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2861" *)
  wire or_tmp_216;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2862" *)
  wire or_tmp_235;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2863" *)
  wire or_tmp_252;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2864" *)
  wire or_tmp_256;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2838" *)
  wire or_tmp_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2839" *)
  wire or_tmp_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2868" *)
  wire or_tmp_291;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2869" *)
  wire or_tmp_296;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2870" *)
  wire or_tmp_315;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2871" *)
  wire or_tmp_332;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2872" *)
  wire or_tmp_336;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2876" *)
  wire or_tmp_371;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2877" *)
  wire or_tmp_376;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2879" *)
  wire or_tmp_395;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2841" *)
  wire or_tmp_40;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2880" *)
  wire or_tmp_411;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2881" *)
  wire or_tmp_415;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2843" *)
  wire or_tmp_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2885" *)
  wire or_tmp_461;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2844" *)
  wire or_tmp_51;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2892" *)
  wire or_tmp_517;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2945" *)
  wire or_tmp_587;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2946" *)
  wire or_tmp_588;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2845" *)
  wire or_tmp_59;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2947" *)
  wire or_tmp_591;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2846" *)
  wire or_tmp_75;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:2847" *)
  wire or_tmp_91;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3255" *)
  reg reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:3278" *)
  reg reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign FpMul_8U_23U_else_2_else_acc_nl = else_MulOp_data_0_lpi_1_dfm_2_30_0_1[30:23] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4565" *) 8'b10000001;
  assign FpMul_8U_23U_p_expo_1_sva_1_mx0w0 = FpMul_8U_23U_else_2_else_acc_nl + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4568" *) MulIn_data_sva_132[30:23];
  assign FpMul_8U_23U_else_2_else_acc_2_nl = else_MulOp_data_1_lpi_1_dfm_2_30_0_1[30:23] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4593" *) 8'b10000001;
  assign FpMul_8U_23U_p_expo_2_sva_1_mx0w0 = FpMul_8U_23U_else_2_else_acc_2_nl + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4596" *) MulIn_data_sva_132[62:55];
  assign FpMul_8U_23U_else_2_else_acc_3_nl = else_MulOp_data_2_lpi_1_dfm_2_30_0_1[30:23] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4621" *) 8'b10000001;
  assign FpMul_8U_23U_p_expo_3_sva_1_mx0w0 = FpMul_8U_23U_else_2_else_acc_3_nl + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4624" *) MulIn_data_sva_132[94:87];
  assign FpMul_8U_23U_else_2_else_acc_4_nl = else_MulOp_data_3_lpi_1_dfm_2_30_0_1[30:23] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4649" *) 8'b10000001;
  assign FpMul_8U_23U_p_expo_sva_1_mx0w0 = FpMul_8U_23U_else_2_else_acc_4_nl + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4652" *) MulIn_data_sva_132[126:119];
  assign mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl = MulIn_data_sva_1[30:23] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4708" *) else_MulOp_data_0_lpi_1_dfm_mx0_30_0[30:23];
  assign mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl = mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl[8:1] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4711" *) 9'b101000001;
  assign mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl = MulIn_data_sva_1[62:55] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4724" *) else_MulOp_data_1_lpi_1_dfm_mx0_30_0[30:23];
  assign mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl = mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl[8:1] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4727" *) 9'b101000001;
  assign mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl = MulIn_data_sva_1[94:87] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4740" *) else_MulOp_data_2_lpi_1_dfm_mx0_30_0[30:23];
  assign mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl = mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl[8:1] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4743" *) 9'b101000001;
  assign mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl = MulIn_data_sva_1[126:119] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4756" *) else_MulOp_data_3_lpi_1_dfm_mx0_30_0[30:23];
  assign mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl = mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl[8:1] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4759" *) 9'b101000001;
  assign mul_mul_1_FpMantRNE_48U_24U_else_acc_nl = else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4773" *) FpMantRNE_48U_24U_else_carry_1_sva_2;
  assign mul_mul_2_FpMantRNE_48U_24U_else_acc_nl = else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4794" *) FpMantRNE_48U_24U_else_carry_2_sva_2;
  assign mul_mul_3_FpMantRNE_48U_24U_else_acc_nl = else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4814" *) FpMantRNE_48U_24U_else_carry_3_sva_2;
  assign mul_mul_4_FpMantRNE_48U_24U_else_acc_nl = else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4834" *) FpMantRNE_48U_24U_else_carry_sva_2;
  assign mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl = FpMul_8U_23U_p_expo_1_sva_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4858" *) 1'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1 = FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4864" *) 1'b1;
  assign mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl = FpMul_8U_23U_p_expo_2_sva_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4880" *) 1'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1 = FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4886" *) 1'b1;
  assign mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl = FpMul_8U_23U_p_expo_3_sva_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4898" *) 1'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1 = FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4904" *) 1'b1;
  assign mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl = FpMul_8U_23U_p_expo_sva_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4916" *) 1'b1;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1 = FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4922" *) 1'b1;
  assign FpMul_8U_23U_oelse_1_acc_nl = else_MulOp_data_0_lpi_1_dfm_mx0_30_0[30:23] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4934" *) 9'b110000001;
  assign mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl = { FpMul_8U_23U_oelse_1_acc_nl[8], FpMul_8U_23U_oelse_1_acc_nl } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4937" *) MulIn_data_sva_1[30:23];
  assign FpMul_8U_23U_oelse_1_acc_1_nl = else_MulOp_data_1_lpi_1_dfm_mx0_30_0[30:23] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4945" *) 9'b110000001;
  assign mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl = { FpMul_8U_23U_oelse_1_acc_1_nl[8], FpMul_8U_23U_oelse_1_acc_1_nl } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4948" *) MulIn_data_sva_1[62:55];
  assign FpMul_8U_23U_oelse_1_acc_2_nl = else_MulOp_data_2_lpi_1_dfm_mx0_30_0[30:23] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4956" *) 9'b110000001;
  assign mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl = { FpMul_8U_23U_oelse_1_acc_2_nl[8], FpMul_8U_23U_oelse_1_acc_2_nl } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4959" *) MulIn_data_sva_1[94:87];
  assign FpMul_8U_23U_oelse_1_acc_3_nl = else_MulOp_data_3_lpi_1_dfm_mx0_30_0[30:23] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4967" *) 9'b110000001;
  assign mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl = { FpMul_8U_23U_oelse_1_acc_3_nl[8], FpMul_8U_23U_oelse_1_acc_3_nl } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4970" *) MulIn_data_sva_1[126:119];
  assign IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva = { IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1086], IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1086:1023] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5500" *) mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  assign IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva = { IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1086], IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1086:1023] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6016" *) mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  assign IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva = { IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1086], IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1086:1023] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6532" *) mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  assign IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva = { IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1086], IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1086:1023] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7048" *) mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_and_nl;
  assign mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = { 1'b1, FpMul_8U_23U_p_expo_1_sva_1_mx0w0[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7051" *) 1'b1;
  assign mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = { 1'b1, FpMul_8U_23U_p_expo_2_sva_1_mx0w0[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7061" *) 1'b1;
  assign mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = { 1'b1, FpMul_8U_23U_p_expo_3_sva_1_mx0w0[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7071" *) 1'b1;
  assign mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl = { 1'b1, FpMul_8U_23U_p_expo_sva_1_mx0w0[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7081" *) 1'b1;
  assign _00374_ = mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *) { asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160 };
  assign _00375_ = mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *) { asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168 };
  assign _00376_ = mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *) { asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164 };
  assign _00377_ = mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *) { asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156 };
  assign _00378_ = else_MulOp_data_slc_else_MulOp_data_0_30_23_5_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *) { and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51 };
  assign _00379_ = else_MulOp_data_slc_else_MulOp_data_1_30_23_5_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *) { and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58 };
  assign _00380_ = else_MulOp_data_slc_else_MulOp_data_2_30_23_5_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *) { and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64 };
  assign _00381_ = else_MulOp_data_slc_else_MulOp_data_3_30_23_5_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10003" *) { and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70 };
  assign _00382_ = MulIn_data_sva_133[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) { or_839_nl, or_839_nl, or_839_nl, or_839_nl, or_839_nl, or_839_nl, or_839_nl, or_839_nl };
  assign _00383_ = MulIn_data_sva_133[62:55] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) { or_838_nl, or_838_nl, or_838_nl, or_838_nl, or_838_nl, or_838_nl, or_838_nl, or_838_nl };
  assign _00384_ = MulIn_data_sva_133[94:87] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) { or_837_nl, or_837_nl, or_837_nl, or_837_nl, or_837_nl, or_837_nl, or_837_nl, or_837_nl };
  assign _00385_ = MulIn_data_sva_133[126:119] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) { or_836_nl, or_836_nl, or_836_nl, or_836_nl, or_836_nl, or_836_nl, or_836_nl, or_836_nl };
  assign _00386_ = else_MulOp_data_0_lpi_1_dfm_2_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) { and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50 };
  assign _00387_ = else_MulOp_data_1_lpi_1_dfm_2_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) { and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57 };
  assign _00388_ = else_MulOp_data_2_lpi_1_dfm_2_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) { and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63 };
  assign _00389_ = else_MulOp_data_3_lpi_1_dfm_2_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) { and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69 };
  assign _00390_ = FpMul_8U_23U_p_expo_1_sva_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) { and_359_nl, and_359_nl, and_359_nl, and_359_nl, and_359_nl, and_359_nl, and_359_nl, and_359_nl };
  assign _00391_ = FpMul_8U_23U_p_expo_2_sva_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) { and_357_nl, and_357_nl, and_357_nl, and_357_nl, and_357_nl, and_357_nl, and_357_nl, and_357_nl };
  assign _00392_ = FpMul_8U_23U_p_expo_3_sva_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) { and_355_nl, and_355_nl, and_355_nl, and_355_nl, and_355_nl, and_355_nl, and_355_nl, and_355_nl };
  assign _00393_ = FpMul_8U_23U_p_expo_sva_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) { and_353_nl, and_353_nl, and_353_nl, and_353_nl, and_353_nl, and_353_nl, and_353_nl, and_353_nl };
  assign _00394_ = FpMul_8U_23U_p_expo_1_sva_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) { and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48 };
  assign _00395_ = FpMul_8U_23U_p_expo_2_sva_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) { and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55 };
  assign _00396_ = FpMul_8U_23U_p_expo_3_sva_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) { and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61 };
  assign _00397_ = FpMul_8U_23U_p_expo_sva_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) { and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67 };
  assign _00398_ = FpMul_8U_23U_FpMul_8U_23U_and_15_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) { and_358_nl, and_358_nl, and_358_nl, and_358_nl, and_358_nl, and_358_nl, and_358_nl, and_358_nl };
  assign _00399_ = FpMul_8U_23U_FpMul_8U_23U_and_16_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) { and_356_nl, and_356_nl, and_356_nl, and_356_nl, and_356_nl, and_356_nl, and_356_nl, and_356_nl };
  assign _00400_ = FpMul_8U_23U_FpMul_8U_23U_and_17_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) { and_354_nl, and_354_nl, and_354_nl, and_354_nl, and_354_nl, and_354_nl, and_354_nl, and_354_nl };
  assign _00401_ = FpMul_8U_23U_FpMul_8U_23U_and_18_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) { and_352_nl, and_352_nl, and_352_nl, and_352_nl, and_352_nl, and_352_nl, and_352_nl, and_352_nl };
  assign _00402_ = FpMul_8U_23U_p_expo_1_sva_1_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) { and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46 };
  assign _00403_ = FpMul_8U_23U_p_expo_2_sva_1_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) { and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54 };
  assign _00404_ = FpMul_8U_23U_p_expo_3_sva_1_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) { and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60 };
  assign _00405_ = FpMul_8U_23U_p_expo_sva_1_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) { and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66 };
  assign _00406_ = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4344" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _00407_ = _00406_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4344" *) or_74_cse;
  assign chn_mul_out_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4344" *) _01023_;
  assign chn_mul_out_and_1_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4345" *) _00753_;
  assign _00408_ = _00754_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4347" *) mul_mul_mul_mul_nor_m1c;
  assign mul_mul_and_m1c = _00408_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4347" *) _00755_;
  assign _00409_ = _00756_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4349" *) mul_mul_mul_mul_nor_2_m1c;
  assign mul_mul_and_17_m1c = _00409_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4349" *) _00755_;
  assign _00410_ = _00757_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4351" *) mul_mul_mul_mul_nor_4_m1c;
  assign mul_mul_and_19_m1c = _00410_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4351" *) _00755_;
  assign _00411_ = _00758_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4353" *) mul_mul_mul_mul_nor_6_m1c;
  assign mul_mul_and_21_m1c = _00411_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4353" *) _00755_;
  assign MulIn_data_and_1_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4354" *) and_18_tmp;
  assign else_MulOp_data_and_8_cse = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4356" *) _00759_;
  assign _00412_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4359" *) IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse;
  assign FpMul_8U_23U_oelse_1_and_4_cse = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4359" *) _00759_;
  assign else_MulOp_data_and_9_cse = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4360" *) _00760_;
  assign FpMul_8U_23U_oelse_1_and_5_cse = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4362" *) _00760_;
  assign else_MulOp_data_and_10_cse = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4363" *) _00761_;
  assign FpMul_8U_23U_oelse_1_and_6_cse = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4365" *) _00761_;
  assign else_MulOp_data_and_11_cse = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4366" *) _00762_;
  assign FpMul_8U_23U_oelse_1_and_7_cse = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4368" *) _00762_;
  assign mul_mul_aelse_and_cse = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4369" *) _00763_;
  assign _00413_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4371" *) _00764_;
  assign MulIn_data_and_2_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4371" *) mux_26_nl;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_8_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4378" *) mux_27_nl;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_9_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4384" *) mux_29_nl;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_10_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4390" *) mux_31_nl;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_11_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4396" *) mux_33_nl;
  assign _00414_ = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4405" *) main_stage_v_2;
  assign IsNaN_8U_23U_1_aelse_and_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4406" *) not_tmp_54;
  assign _00415_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4410" *) FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse;
  assign FpMantRNE_48U_24U_else_and_cse = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4410" *) not_tmp_55;
  assign IsNaN_8U_23U_aelse_and_17_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4414" *) _00770_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_13_cse = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4416" *) not_tmp_54;
  assign _00416_ = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4424" *) main_stage_v_2;
  assign IsNaN_8U_23U_1_aelse_and_1_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4425" *) not_tmp_81;
  assign FpMantRNE_48U_24U_else_and_9_cse = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4429" *) not_tmp_82;
  assign IsNaN_8U_23U_aelse_and_19_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4433" *) _00774_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_16_cse = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4435" *) not_tmp_81;
  assign _00417_ = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4443" *) main_stage_v_2;
  assign IsNaN_8U_23U_1_aelse_and_2_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4444" *) not_tmp_106;
  assign FpMantRNE_48U_24U_else_and_11_cse = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4448" *) not_tmp_107;
  assign IsNaN_8U_23U_aelse_and_21_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4452" *) _00778_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_19_cse = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4454" *) not_tmp_106;
  assign IsNaN_8U_23U_1_aelse_and_3_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4463" *) not_tmp_129;
  assign FpMantRNE_48U_24U_else_and_13_cse = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4467" *) not_tmp_130;
  assign IsNaN_8U_23U_aelse_and_23_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4471" *) _00782_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_22_cse = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4473" *) not_tmp_129;
  assign mul_mul_aelse_and_12_cse = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4474" *) _00783_;
  assign MulIn_data_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4475" *) _00785_;
  assign IsNaN_8U_23U_aelse_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4476" *) _00786_;
  assign _00418_ = IsNaN_8U_23U_aelse_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4481" *) IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_3_cse;
  assign IsNaN_8U_23U_aelse_and_24_cse = _00418_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4481" *) _00787_;
  assign IsNaN_8U_23U_aelse_and_25_cse = _00418_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4485" *) _00788_;
  assign IsNaN_8U_23U_aelse_and_26_cse = _00418_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4489" *) _00789_;
  assign IsNaN_8U_23U_aelse_and_27_cse = _00418_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4493" *) _00790_;
  assign _00419_ = IsNaN_8U_23U_aelse_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4494" *) and_20_tmp;
  assign mul_mul_aelse_and_19_cse = _00419_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4495" *) _00791_;
  assign FpMul_8U_23U_p_expo_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4497" *) _00792_;
  assign else_MulOp_data_and_1_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4498" *) _00793_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4500" *) _00794_;
  assign FpMul_8U_23U_p_expo_and_1_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4501" *) _00795_;
  assign else_MulOp_data_and_3_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4502" *) _00796_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_2_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4504" *) _00797_;
  assign FpMul_8U_23U_p_expo_and_2_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4505" *) _00798_;
  assign else_MulOp_data_and_5_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4506" *) _00799_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_4_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4508" *) _00800_;
  assign FpMul_8U_23U_p_expo_and_3_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4509" *) _00801_;
  assign else_MulOp_data_and_7_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4510" *) _00802_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_6_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4512" *) _00803_;
  assign and_136_m1c = and_18_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4513" *) _00804_;
  assign and_135_rgt = and_18_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4514" *) IsNaN_8U_23U_land_1_lpi_1_dfm_4;
  assign mul_mul_if_and_6_rgt = _00805_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4515" *) and_136_m1c;
  assign mul_mul_if_and_7_rgt = IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4516" *) and_136_m1c;
  assign and_138_m1c = and_18_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4517" *) _00806_;
  assign and_137_rgt = and_18_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4518" *) IsNaN_8U_23U_land_2_lpi_1_dfm_4;
  assign mul_mul_if_and_4_rgt = _00807_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4519" *) and_138_m1c;
  assign mul_mul_if_and_5_rgt = IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4520" *) and_138_m1c;
  assign and_140_m1c = and_18_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4521" *) _00808_;
  assign and_139_rgt = and_18_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4522" *) IsNaN_8U_23U_land_3_lpi_1_dfm_4;
  assign mul_mul_if_and_2_rgt = _00809_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4523" *) and_140_m1c;
  assign mul_mul_if_and_3_rgt = IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4524" *) and_140_m1c;
  assign and_142_m1c = and_18_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4525" *) _00810_;
  assign and_141_rgt = and_18_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4526" *) IsNaN_8U_23U_land_lpi_1_dfm_4;
  assign mul_mul_if_and_rgt = _00811_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4527" *) and_142_m1c;
  assign mul_mul_if_and_1_rgt = IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4528" *) and_142_m1c;
  assign and_146_rgt = _01068_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4532" *) and_18_tmp;
  assign and_150_rgt = _01069_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4536" *) and_18_tmp;
  assign and_154_rgt = _01070_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4540" *) and_18_tmp;
  assign and_158_rgt = _01072_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4544" *) and_18_tmp;
  assign _00420_ = cfg_mul_prelu_rsci_d & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *) _00816_;
  assign IsNaN_8U_23U_aelse_and_4_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *) _00817_;
  assign _00421_ = cfg_mul_prelu_rsci_d & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *) _00818_;
  assign IsNaN_8U_23U_aelse_and_5_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *) _00819_;
  assign _00422_ = cfg_mul_prelu_rsci_d & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *) _00820_;
  assign IsNaN_8U_23U_aelse_and_6_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *) _00821_;
  assign _00423_ = cfg_mul_prelu_rsci_d & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *) _00822_;
  assign IsNaN_8U_23U_aelse_and_7_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *) _00823_;
  assign _00424_ = mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4571" *) mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign mul_mul_1_FpMantRNE_48U_24U_else_and_tmp = FpMantRNE_48U_24U_else_carry_1_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4573" *) _00708_;
  assign _00425_ = FpMul_8U_23U_p_mant_p1_1_sva_mx1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4575" *) FpMul_8U_23U_p_mant_p1_1_sva_mx1[47];
  assign FpMantRNE_48U_24U_else_carry_1_sva_mx0w0 = FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4587" *) _01107_;
  assign FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0 = _01108_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4589" *) mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign _00426_ = mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4599" *) mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign mul_mul_2_FpMantRNE_48U_24U_else_and_tmp = FpMantRNE_48U_24U_else_carry_2_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4601" *) _00710_;
  assign _00427_ = FpMul_8U_23U_p_mant_p1_2_sva_mx1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4603" *) FpMul_8U_23U_p_mant_p1_2_sva_mx1[47];
  assign FpMantRNE_48U_24U_else_carry_2_sva_mx0w0 = FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4615" *) _01131_;
  assign FpMul_8U_23U_FpMul_8U_23U_and_12_itm_mx0w0 = _01132_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4617" *) mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign _00428_ = mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4627" *) mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign mul_mul_3_FpMantRNE_48U_24U_else_and_tmp = FpMantRNE_48U_24U_else_carry_3_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4629" *) _00712_;
  assign _00429_ = FpMul_8U_23U_p_mant_p1_3_sva_mx1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4631" *) FpMul_8U_23U_p_mant_p1_3_sva_mx1[47];
  assign FpMantRNE_48U_24U_else_carry_3_sva_mx0w0 = FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4643" *) _01155_;
  assign FpMul_8U_23U_FpMul_8U_23U_and_13_itm_mx0w0 = _01156_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4645" *) mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign _00430_ = mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4655" *) mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign mul_mul_4_FpMantRNE_48U_24U_else_and_tmp = FpMantRNE_48U_24U_else_carry_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4657" *) _00714_;
  assign _00431_ = FpMul_8U_23U_p_mant_p1_sva_mx1[0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4659" *) FpMul_8U_23U_p_mant_p1_sva_mx1[47];
  assign FpMantRNE_48U_24U_else_carry_sva_mx0w0 = FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4671" *) _01179_;
  assign FpMul_8U_23U_FpMul_8U_23U_and_14_itm_mx0w0 = _01180_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4673" *) mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign FpMul_8U_23U_p_mant_p1_and_7_nl = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4701" *) _00829_;
  assign FpMul_8U_23U_p_mant_p1_and_6_nl = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4717" *) _00832_;
  assign FpMul_8U_23U_p_mant_p1_and_5_nl = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4733" *) _00835_;
  assign FpMul_8U_23U_p_mant_p1_and_4_nl = mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4749" *) _00838_;
  assign FpMul_8U_23U_and_1_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4784" *) _00754_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_64_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4791" *) mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign FpMul_8U_23U_and_3_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4805" *) _00756_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_64_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4812" *) mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign FpMul_8U_23U_and_5_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4825" *) _00757_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_64_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4832" *) mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign FpMul_8U_23U_and_7_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4845" *) _00758_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_64_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4852" *) mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign _00432_ = _00011_[22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4869" *) mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2;
  assign _00433_ = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4871" *) mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl = _00433_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4871" *) or_tmp_133;
  assign _00434_ = _00014_[22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4889" *) mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2;
  assign _00435_ = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4891" *) mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl = _00435_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4891" *) _00846_;
  assign _00436_ = _00017_[22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4907" *) mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2;
  assign _00437_ = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4909" *) mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl = _00437_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4909" *) _00848_;
  assign _00438_ = _00020_[22] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4925" *) mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2;
  assign _00439_ = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4927" *) mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl = _00439_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4927" *) _00850_;
  assign _00440_ = chn_mul_in_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4977" *) or_11_cse;
  assign _00441_ = _00440_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4977" *) or_12_cse;
  assign _00442_ = _00441_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4977" *) or_13_cse;
  assign _00443_ = _00442_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4978" *) or_14_cse;
  assign _00444_ = _00443_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4978" *) or_15_cse;
  assign _00445_ = _00444_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4978" *) or_16_cse;
  assign and_20_tmp = _00445_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4978" *) or_74_cse;
  assign _00446_ = cfg_mul_src_1_sva_st_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4980" *) _00763_;
  assign _00447_ = _00446_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4980" *) main_stage_v_1;
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_and_nl = IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1022] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5498" *) _02224_;
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_and_nl = IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1022] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6014" *) _03246_;
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_and_nl = IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1022] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6530" *) _04268_;
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_and_nl = IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1022] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7046" *) _05290_;
  assign _00448_ = mul_mul_else_unequal_tmp_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7088" *) _00858_;
  assign asn_156 = _00448_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7089" *) _00755_;
  assign _00449_ = mul_mul_else_unequal_tmp_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7091" *) _00859_;
  assign asn_160 = _00449_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7092" *) _00755_;
  assign _00450_ = mul_mul_else_unequal_tmp_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7094" *) _00860_;
  assign asn_164 = _00450_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7095" *) _00755_;
  assign _00451_ = mul_mul_else_unequal_tmp_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7097" *) _00861_;
  assign asn_168 = _00451_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7098" *) _00755_;
  assign _00452_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7100" *) or_11_cse;
  assign _00453_ = _00452_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7100" *) or_12_cse;
  assign _00454_ = _00453_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7100" *) or_13_cse;
  assign _00455_ = _00454_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7101" *) or_14_cse;
  assign _00456_ = _00455_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7101" *) or_15_cse;
  assign _00457_ = _00456_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7101" *) or_16_cse;
  assign and_18_tmp = _00457_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7101" *) or_74_cse;
  assign _00458_ = mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7180" *) FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_3;
  assign _00459_ = mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7271" *) main_stage_v_2;
  assign and_dcpl_3 = and_20_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7298" *) and_dcpl_37;
  assign and_dcpl_6 = or_27_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7300" *) and_20_tmp;
  assign and_tmp_5 = FpMul_8U_23U_FpMul_8U_23U_and_14_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7305" *) or_tmp_411;
  assign _00460_ = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7306" *) _00755_;
  assign and_dcpl_22 = _00460_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7306" *) or_74_cse;
  assign and_dcpl_23 = _00869_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7307" *) reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign and_dcpl_24 = or_74_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7308" *) main_stage_v_3;
  assign _00461_ = _00752_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7309" *) chn_mul_out_rsci_bawt;
  assign and_dcpl_26 = _00461_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7309" *) reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign and_dcpl_27 = _00791_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7310" *) and_20_tmp;
  assign and_dcpl_30 = _00446_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7313" *) and_18_tmp;
  assign and_dcpl_38 = and_dcpl_37 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7316" *) and_18_tmp;
  assign and_dcpl_39 = or_27_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7317" *) and_18_tmp;
  assign and_dcpl_45 = or_74_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7318" *) _00870_;
  assign _00462_ = and_dcpl_45 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7319" *) cfg_precision[1];
  assign and_dcpl_46 = _00462_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7319" *) _00871_;
  assign and_dcpl_47 = or_74_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7320" *) or_27_cse;
  assign and_dcpl_48 = and_dcpl_47 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7321" *) _00871_;
  assign and_dcpl_50 = _00462_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7322" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign and_dcpl_51 = and_dcpl_47 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7323" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign and_dcpl_52 = or_74_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7324" *) and_dcpl_37;
  assign and_dcpl_54 = _00462_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7325" *) _00872_;
  assign and_dcpl_55 = and_dcpl_47 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7326" *) _00872_;
  assign and_dcpl_57 = _00462_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7327" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign and_dcpl_58 = and_dcpl_47 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7328" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign and_dcpl_60 = _00462_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7329" *) _00873_;
  assign and_dcpl_61 = and_dcpl_47 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7330" *) _00873_;
  assign and_dcpl_63 = _00462_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7331" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign and_dcpl_64 = and_dcpl_47 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7332" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign and_dcpl_66 = _00462_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7333" *) _00874_;
  assign and_dcpl_67 = and_dcpl_47 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7334" *) _00874_;
  assign and_dcpl_69 = _00462_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7335" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign and_dcpl_70 = and_dcpl_47 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7336" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _00463_ = cfg_precision[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7359" *) and_18_tmp;
  assign or_tmp_587 = and_20_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7366" *) fsm_output[1];
  assign _00464_ = and_dcpl_27 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7367" *) cfg_mul_src_rsci_d;
  assign or_tmp_588 = _00464_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7367" *) fsm_output[1];
  assign or_tmp_591 = and_18_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7368" *) fsm_output[1];
  assign chn_mul_op_rsci_ld_core_psct_mx0c1 = and_dcpl_30 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7370" *) _05463_;
  assign _00465_ = or_74_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7371" *) main_stage_v_2;
  assign main_stage_v_2_mx0c1 = _00465_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7371" *) _00812_;
  assign _00466_ = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7372" *) _00766_;
  assign main_stage_v_3_mx0c1 = _00466_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7372" *) or_74_cse;
  assign _00467_ = _00784_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7373" *) and_18_tmp;
  assign main_stage_v_1_mx0c1 = _00467_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7373" *) fsm_output[1];
  assign _00468_ = cfg_mul_bypass_rsci_d & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7374" *) and_20_tmp;
  assign cfg_mul_src_1_sva_st_1_mx0c1 = _00468_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7374" *) fsm_output[1];
  assign chn_mul_out_rsci_oswt_unreg = chn_mul_out_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7377" *) reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign _00469_ = _00784_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7387" *) fsm_output[1];
  assign _00470_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7397" *) chn_mul_in_rsci_ld_core_psct_mx0c0;
  assign _00471_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7473" *) _05464_;
  assign _00472_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7481" *) _05465_;
  assign _00473_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7489" *) _05466_;
  assign _00474_ = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7497" *) not_tmp_2;
  assign _00475_ = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7532" *) not_tmp_2;
  assign _00476_ = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7553" *) _00881_;
  assign _00477_ = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7575" *) not_tmp_8;
  assign _00478_ = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7584" *) not_tmp_8;
  assign _00479_ = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7605" *) _00882_;
  assign _00480_ = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7627" *) not_tmp_12;
  assign _00481_ = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7636" *) not_tmp_12;
  assign _00482_ = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7657" *) _00883_;
  assign _00483_ = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7679" *) not_tmp_15;
  assign _00484_ = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7688" *) not_tmp_15;
  assign _00485_ = _00412_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7709" *) _00884_;
  assign _00486_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7745" *) _05467_;
  assign _00487_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7820" *) FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_3_cse;
  assign _00488_ = _00487_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7821" *) mux_42_nl;
  assign _00489_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7834" *) mux_44_nl;
  assign _00490_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7846" *) mux_49_nl;
  assign _00491_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7856" *) mux_50_nl;
  assign _00492_ = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7866" *) _00886_;
  assign _00493_ = _00487_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7897" *) mux_63_nl;
  assign _00494_ = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7918" *) not_tmp_55;
  assign _00495_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7927" *) _00770_;
  assign _00496_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7936" *) mux_66_nl;
  assign _00497_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7957" *) FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_2_cse;
  assign _00498_ = _00497_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7958" *) mux_74_nl;
  assign _00499_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7971" *) mux_76_nl;
  assign _00500_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7983" *) mux_81_nl;
  assign _00501_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7993" *) mux_82_nl;
  assign _00502_ = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8003" *) _00887_;
  assign _00503_ = _00497_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8034" *) mux_93_nl;
  assign _00504_ = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8055" *) not_tmp_82;
  assign _00505_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8064" *) _00774_;
  assign _00506_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8073" *) mux_97_nl;
  assign _00507_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8094" *) FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_1_cse;
  assign _00508_ = _00507_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8095" *) mux_105_nl;
  assign _00509_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8108" *) mux_107_nl;
  assign _00510_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8120" *) mux_112_nl;
  assign _00511_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8130" *) mux_113_nl;
  assign _00512_ = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8140" *) _00888_;
  assign _00513_ = _00507_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8171" *) mux_124_nl;
  assign _00514_ = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8192" *) not_tmp_107;
  assign _00515_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8201" *) _00778_;
  assign _00516_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8210" *) mux_128_nl;
  assign _00517_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8231" *) FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_cse;
  assign _00518_ = _00517_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8232" *) mux_136_nl;
  assign _00519_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8245" *) mux_138_nl;
  assign _00520_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8257" *) mux_143_nl;
  assign _00521_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8267" *) _00889_;
  assign _00522_ = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8277" *) _00890_;
  assign _00523_ = _00517_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8308" *) mux_156_nl;
  assign _00524_ = _00413_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8329" *) not_tmp_130;
  assign _00525_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8338" *) _00782_;
  assign _00526_ = _00415_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8347" *) mux_159_nl;
  assign _00527_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8382" *) _05468_;
  assign _00528_ = _00419_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8431" *) _00892_;
  assign _00529_ = _00419_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8439" *) _00893_;
  assign _00530_ = and_dcpl_27 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8497" *) fsm_output[1];
  assign _00531_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8498" *) _05470_;
  assign _00532_ = FpMul_8U_23U_p_expo_and_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8508" *) mux_185_nl;
  assign _00533_ = else_MulOp_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8518" *) mux_187_nl;
  assign _00534_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8540" *) _00894_;
  assign _00535_ = FpMul_8U_23U_p_expo_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8573" *) mux_189_nl;
  assign _00536_ = else_MulOp_data_and_3_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8583" *) mux_191_nl;
  assign _00537_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8605" *) _00895_;
  assign _00538_ = FpMul_8U_23U_p_expo_and_2_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8638" *) mux_193_nl;
  assign _00539_ = else_MulOp_data_and_5_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8648" *) mux_195_nl;
  assign _00540_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8670" *) _00896_;
  assign _00541_ = FpMul_8U_23U_p_expo_and_3_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8703" *) mux_197_nl;
  assign _00542_ = else_MulOp_data_and_7_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8713" *) mux_201_nl;
  assign _00543_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8735" *) _00897_;
  assign _00544_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8767" *) mux_203_nl;
  assign _00545_ = FpMul_8U_23U_oelse_1_mux_20_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8768" *) _00898_;
  assign _00546_ = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8776" *) _00899_;
  assign _00547_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8785" *) _05481_;
  assign _00548_ = _00547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8785" *) mux_207_nl;
  assign _00549_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8795" *) mux_209_nl;
  assign _00550_ = FpMul_8U_23U_oelse_1_mux_21_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8796" *) _00898_;
  assign _00551_ = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8804" *) _00900_;
  assign _00552_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8813" *) _05485_;
  assign _00553_ = _00552_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8813" *) mux_213_nl;
  assign _00554_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8823" *) mux_215_nl;
  assign _00555_ = FpMul_8U_23U_oelse_1_mux_22_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8824" *) _00898_;
  assign _00556_ = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8832" *) _00901_;
  assign _00557_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8841" *) _05489_;
  assign _00558_ = _00557_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8841" *) mux_219_nl;
  assign _00559_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8851" *) mux_221_nl;
  assign _00560_ = FpMul_8U_23U_oelse_1_mux_23_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8852" *) _00898_;
  assign _00561_ = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8860" *) _00902_;
  assign _00562_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8869" *) _05493_;
  assign _00563_ = _00562_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8869" *) mux_225_nl;
  assign _00564_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8880" *) _00903_;
  assign _00565_ = _00564_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8881" *) mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign _00566_ = nor_118_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8890" *) and_dcpl_38;
  assign _00567_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8890" *) _05497_;
  assign _00568_ = _00567_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8891" *) _00759_;
  assign _00569_ = mul_mul_land_2_lpi_1_dfm_st_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8902" *) mul_mul_land_lpi_1_dfm_st_1;
  assign _00570_ = _00569_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8902" *) mul_mul_land_1_lpi_1_dfm_st_1;
  assign _00571_ = _00570_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8902" *) mul_mul_land_3_lpi_1_dfm_st_1;
  assign _00572_ = MulIn_data_and_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8903" *) _00904_;
  assign _00573_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8911" *) _00905_;
  assign _00574_ = _00573_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8912" *) mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign _00575_ = nor_117_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8921" *) and_dcpl_38;
  assign _00576_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8921" *) _05501_;
  assign _00577_ = _00576_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8922" *) _00760_;
  assign _00578_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8932" *) _00906_;
  assign _00579_ = _00578_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8933" *) mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign _00580_ = nor_116_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8942" *) and_dcpl_38;
  assign _00581_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8942" *) _05504_;
  assign _00582_ = _00581_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8943" *) _00761_;
  assign _00583_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8954" *) _00907_;
  assign _00584_ = _00583_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8955" *) mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign _00585_ = nor_115_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8964" *) and_dcpl_38;
  assign _00586_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8964" *) _05507_;
  assign _00587_ = _00586_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8965" *) _00762_;
  assign _00588_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8975" *) _00908_;
  assign _00589_ = _00588_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8975" *) _00909_;
  assign _00590_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8983" *) _00910_;
  assign _00591_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8991" *) _00911_;
  assign _00592_ = _00591_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8991" *) _00912_;
  assign _00593_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8999" *) _00913_;
  assign _00594_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9007" *) _00914_;
  assign _00595_ = _00594_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9007" *) _00915_;
  assign _00596_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9015" *) _00916_;
  assign _00597_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9023" *) _00917_;
  assign _00598_ = _00597_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9023" *) _00918_;
  assign _00599_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9031" *) _00919_;
  assign _00600_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9079" *) _00920_;
  assign _00601_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9089" *) _00921_;
  assign _00602_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9098" *) _00922_;
  assign _00603_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9108" *) _00923_;
  assign _00604_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9117" *) _00924_;
  assign _00605_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9127" *) _00925_;
  assign _00606_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9136" *) _00926_;
  assign _00607_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9146" *) _00927_;
  assign _00608_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9155" *) _00928_;
  assign and_358_nl = _00937_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9233" *) mul_mul_and_m1c;
  assign and_359_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9234" *) mul_mul_and_m1c;
  assign _00609_ = IsNaN_8U_23U_land_1_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9235" *) mul_mul_mul_mul_nor_m1c;
  assign _00610_ = _00609_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9236" *) _00755_;
  assign and_356_nl = _00938_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9251" *) mul_mul_and_17_m1c;
  assign and_357_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9252" *) mul_mul_and_17_m1c;
  assign _00611_ = IsNaN_8U_23U_land_2_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9254" *) mul_mul_mul_mul_nor_2_m1c;
  assign _00612_ = _00611_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9254" *) _00755_;
  assign and_354_nl = _00939_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9269" *) mul_mul_and_19_m1c;
  assign and_355_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9270" *) mul_mul_and_19_m1c;
  assign _00613_ = IsNaN_8U_23U_land_3_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9272" *) mul_mul_mul_mul_nor_4_m1c;
  assign _00614_ = _00613_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9272" *) _00755_;
  assign and_352_nl = _00940_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9287" *) mul_mul_and_21_m1c;
  assign and_353_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9288" *) mul_mul_and_21_m1c;
  assign _00615_ = IsNaN_8U_23U_land_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9289" *) mul_mul_mul_mul_nor_6_m1c;
  assign _00616_ = _00615_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9290" *) _00755_;
  assign _00617_ = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9331" *) mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign and_344_nl = _00944_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9338" *) mux_39_nl;
  assign _00618_ = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9343" *) mux_40_nl;
  assign _00619_ = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9357" *) mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  assign _00620_ = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9375" *) _05615_;
  assign _00621_ = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9393" *) mux_60_nl;
  assign and_343_nl = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9413" *) mux_64_nl;
  assign _00622_ = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9435" *) mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign _00623_ = mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9444" *) FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_3;
  assign _00624_ = _00623_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9444" *) _00959_;
  assign and_342_nl = _00624_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9444" *) mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign _00625_ = _05675_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9447" *) mux_72_nl;
  assign _00626_ = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9461" *) mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  assign _00627_ = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9497" *) mux_90_nl;
  assign and_340_nl = _00964_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9504" *) mux_92_nl;
  assign and_339_nl = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9518" *) mux_95_nl;
  assign _00628_ = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9540" *) mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign _00629_ = mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9549" *) FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_3;
  assign _00630_ = _00629_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9549" *) _00972_;
  assign and_338_nl = _00630_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9549" *) mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign _00631_ = _05759_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9552" *) mux_103_nl;
  assign _00632_ = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9566" *) mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  assign _00633_ = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9602" *) mux_121_nl;
  assign and_336_nl = _00977_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9609" *) mux_123_nl;
  assign and_335_nl = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9623" *) mux_126_nl;
  assign _00634_ = FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9645" *) mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign _00635_ = mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9654" *) FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_3;
  assign _00636_ = _00635_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9654" *) _00985_;
  assign and_334_nl = _00636_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9654" *) mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign _00637_ = _05842_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9657" *) mux_134_nl;
  assign _00638_ = mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9671" *) mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  assign _00639_ = mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9708" *) mux_153_nl;
  assign and_332_nl = _00990_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9715" *) mux_155_nl;
  assign and_331_nl = mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9729" *) mux_157_nl;
  assign and_39_nl = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9751" *) mux_186_nl;
  assign and_40_nl = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9769" *) mux_190_nl;
  assign and_41_nl = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9787" *) mux_194_nl;
  assign and_328_nl = _01056_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9804" *) mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign _00640_ = _00732_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9813" *) _00716_;
  assign _00641_ = _00734_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9831" *) _00717_;
  assign _00642_ = _00736_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9849" *) _00718_;
  assign _00643_ = _00738_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9867" *) _00719_;
  assign _00644_ = else_MulOp_data_0_lpi_1_dfm_mx1[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9935" *) mul_mul_if_and_7_rgt;
  assign _00645_ = else_MulOp_data_1_lpi_1_dfm_mx1[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9935" *) mul_mul_if_and_5_rgt;
  assign _00646_ = else_MulOp_data_2_lpi_1_dfm_mx1[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9935" *) mul_mul_if_and_3_rgt;
  assign _00647_ = else_MulOp_data_3_lpi_1_dfm_mx1[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9935" *) mul_mul_if_and_1_rgt;
  assign _00648_ = mul_mul_1_FpMul_8U_23U_xor_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *) mul_mul_if_and_6_rgt;
  assign _00649_ = mul_mul_2_FpMul_8U_23U_xor_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *) mul_mul_if_and_4_rgt;
  assign _00650_ = mul_mul_3_FpMul_8U_23U_xor_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *) mul_mul_if_and_2_rgt;
  assign _00651_ = mul_mul_4_FpMul_8U_23U_xor_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *) mul_mul_if_and_rgt;
  assign _00652_ = MulIn_data_sva_1[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *) and_135_rgt;
  assign _00653_ = MulIn_data_sva_1[63] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *) and_137_rgt;
  assign _00654_ = MulIn_data_sva_1[95] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *) and_139_rgt;
  assign _00655_ = MulIn_data_sva_1[127] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *) and_141_rgt;
  assign _00656_ = MulIn_data_sva_133[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9948" *) { asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162, asn_162 };
  assign _00657_ = MulIn_data_sva_133[54:33] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9948" *) { asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170, asn_170 };
  assign _00658_ = MulIn_data_sva_133[86:65] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9948" *) { asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166, asn_166 };
  assign _00659_ = MulIn_data_sva_133[118:97] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9948" *) { asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158, asn_158 };
  assign _00660_ = mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *) { asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160, asn_160 };
  assign _00661_ = mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *) { asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168, asn_168 };
  assign _00662_ = mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *) { asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164, asn_164 };
  assign _00663_ = mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *) { asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156, asn_156 };
  assign _00664_ = FpMul_8U_23U_o_mant_1_lpi_1_dfm_3[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *) { nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl, nor_3_nl };
  assign _00665_ = FpMul_8U_23U_o_mant_2_lpi_1_dfm_3[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *) { nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl, nor_2_nl };
  assign _00666_ = FpMul_8U_23U_o_mant_3_lpi_1_dfm_3[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *) { nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl, nor_1_nl };
  assign _00667_ = FpMul_8U_23U_o_mant_lpi_1_dfm_3[22:1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *) { nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl, nor_6_nl };
  assign _00668_ = MulIn_data_sva_133[22:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9961" *) { IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8, IsNaN_8U_23U_land_1_lpi_1_dfm_8 };
  assign _00669_ = MulIn_data_sva_133[54:32] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9961" *) { IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8, IsNaN_8U_23U_land_2_lpi_1_dfm_8 };
  assign _00670_ = MulIn_data_sva_133[86:64] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9961" *) { IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8, IsNaN_8U_23U_land_3_lpi_1_dfm_8 };
  assign _00671_ = MulIn_data_sva_133[118:96] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9961" *) { IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8, IsNaN_8U_23U_land_lpi_1_dfm_8 };
  assign _00672_ = else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *) { FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl, FpMul_8U_23U_and_1_nl };
  assign _00673_ = else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *) { FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl, FpMul_8U_23U_and_3_nl };
  assign _00674_ = else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *) { FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl, FpMul_8U_23U_and_5_nl };
  assign _00675_ = else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *) { FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl, FpMul_8U_23U_and_7_nl };
  assign _00676_ = FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *) { FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl, FpMul_8U_23U_FpMul_8U_23U_nor_nl };
  assign _00677_ = FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *) { FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl, FpMul_8U_23U_FpMul_8U_23U_nor_1_nl };
  assign _00678_ = FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_6_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *) { FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl, FpMul_8U_23U_FpMul_8U_23U_nor_2_nl };
  assign _00679_ = FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *) { FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl, FpMul_8U_23U_FpMul_8U_23U_nor_3_nl };
  assign _00680_ = mul_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9975" *) { and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48, and_dcpl_48 };
  assign _00681_ = mul_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9975" *) { and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55, and_dcpl_55 };
  assign _00682_ = mul_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9975" *) { and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61, and_dcpl_61 };
  assign _00683_ = mul_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9975" *) { and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67, and_dcpl_67 };
  assign _00684_ = FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[45:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *) { and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46, and_dcpl_46 };
  assign _00685_ = FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[45:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *) { and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54, and_dcpl_54 };
  assign _00686_ = FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[45:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *) { and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60, and_dcpl_60 };
  assign _00687_ = FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[45:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *) { and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66, and_dcpl_66 };
  assign _00688_ = else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *) { and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51, and_dcpl_51 };
  assign _00689_ = else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *) { and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58, and_dcpl_58 };
  assign _00690_ = else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *) { and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64, and_dcpl_64 };
  assign _00691_ = else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *) { and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70, and_dcpl_70 };
  assign _00692_ = else_MulOp_data_0_lpi_1_dfm_2_30_0_1[22:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *) { and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50, and_dcpl_50 };
  assign _00693_ = else_MulOp_data_1_lpi_1_dfm_2_30_0_1[22:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *) { and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57, and_dcpl_57 };
  assign _00694_ = else_MulOp_data_2_lpi_1_dfm_2_30_0_1[22:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *) { and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63, and_dcpl_63 };
  assign _00695_ = else_MulOp_data_3_lpi_1_dfm_2_30_0_1[22:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *) { and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69, and_dcpl_69 };
  assign _00696_ = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9989" *) { FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_1_nl };
  assign _00697_ = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9989" *) { FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_3_nl };
  assign _00698_ = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9989" *) { FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_5_nl };
  assign _00699_ = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9989" *) { FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl, FpMantWidthDec_8U_47U_23U_0U_0U_and_7_nl };
  assign _00700_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *) { FpMul_8U_23U_or_4_nl, FpMul_8U_23U_or_4_nl, FpMul_8U_23U_or_4_nl, FpMul_8U_23U_or_4_nl, FpMul_8U_23U_or_4_nl, FpMul_8U_23U_or_4_nl, FpMul_8U_23U_or_4_nl, FpMul_8U_23U_or_4_nl };
  assign _00701_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *) { FpMul_8U_23U_or_5_nl, FpMul_8U_23U_or_5_nl, FpMul_8U_23U_or_5_nl, FpMul_8U_23U_or_5_nl, FpMul_8U_23U_or_5_nl, FpMul_8U_23U_or_5_nl, FpMul_8U_23U_or_5_nl, FpMul_8U_23U_or_5_nl };
  assign _00702_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *) { FpMul_8U_23U_or_6_nl, FpMul_8U_23U_or_6_nl, FpMul_8U_23U_or_6_nl, FpMul_8U_23U_or_6_nl, FpMul_8U_23U_or_6_nl, FpMul_8U_23U_or_6_nl, FpMul_8U_23U_or_6_nl, FpMul_8U_23U_or_6_nl };
  assign _00703_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *) { FpMul_8U_23U_or_7_nl, FpMul_8U_23U_or_7_nl, FpMul_8U_23U_or_7_nl, FpMul_8U_23U_or_7_nl, FpMul_8U_23U_or_7_nl, FpMul_8U_23U_or_7_nl, FpMul_8U_23U_or_7_nl, FpMul_8U_23U_or_7_nl };
  assign _00704_ = FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *) { FpMul_8U_23U_FpMul_8U_23U_nor_4_nl, FpMul_8U_23U_FpMul_8U_23U_nor_4_nl, FpMul_8U_23U_FpMul_8U_23U_nor_4_nl, FpMul_8U_23U_FpMul_8U_23U_nor_4_nl, FpMul_8U_23U_FpMul_8U_23U_nor_4_nl, FpMul_8U_23U_FpMul_8U_23U_nor_4_nl, FpMul_8U_23U_FpMul_8U_23U_nor_4_nl, FpMul_8U_23U_FpMul_8U_23U_nor_4_nl };
  assign _00705_ = FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *) { nor_267_cse, nor_267_cse, nor_267_cse, nor_267_cse, nor_267_cse, nor_267_cse, nor_267_cse, nor_267_cse };
  assign _00706_ = FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *) { nor_230_cse, nor_230_cse, nor_230_cse, nor_230_cse, nor_230_cse, nor_230_cse, nor_230_cse, nor_230_cse };
  assign _00707_ = FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *) { nor_193_cse, nor_193_cse, nor_193_cse, nor_193_cse, nor_193_cse, nor_193_cse, nor_193_cse, nor_193_cse };
  assign _00708_ = FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[45:23] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4573" *) 23'b11111111111111111111111;
  assign _00709_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva[63:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4590" *) 33'b111111111111111111111111111111111;
  assign _00710_ = FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[45:23] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4601" *) 23'b11111111111111111111111;
  assign _00711_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva[63:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4618" *) 33'b111111111111111111111111111111111;
  assign _00712_ = FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[45:23] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4629" *) 23'b11111111111111111111111;
  assign _00713_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva[63:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4646" *) 33'b111111111111111111111111111111111;
  assign _00714_ = FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[45:23] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4657" *) 23'b11111111111111111111111;
  assign _00715_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva[63:31] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4674" *) 33'b111111111111111111111111111111111;
  assign and_dcpl_37 = cfg_precision == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4792" *) 2'b10;
  assign _00011_[22] = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4862" *) 8'b11111111;
  assign _00014_[22] = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4884" *) 8'b11111111;
  assign _00017_[22] = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4902" *) 8'b11111111;
  assign _00020_[22] = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4920" *) 8'b11111111;
  assign _00716_ = else_mux_tmp_30_23 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9813" *) 8'b11111111;
  assign _00717_ = else_mux_1_tmp_30_23 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9831" *) 8'b11111111;
  assign _00718_ = else_mux_2_tmp_30_23 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9849" *) 8'b11111111;
  assign _00719_ = else_mux_3_tmp_30_23 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9867" *) 8'b11111111;
  assign mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp = { _00830_, MulIn_data_sva_132[22:0] } * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4706" *) { _00831_, else_MulOp_data_0_lpi_1_dfm_2_30_0_1[22:0] };
  assign mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 = $signed(MulIn_data_sva_1[31:0]) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4715" *) $signed(else_MulOp_data_0_lpi_1_dfm_mx1);
  assign mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp = { _00833_, MulIn_data_sva_132[54:32] } * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4722" *) { _00834_, else_MulOp_data_1_lpi_1_dfm_2_30_0_1[22:0] };
  assign mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 = $signed(MulIn_data_sva_1[63:32]) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4731" *) $signed(else_MulOp_data_1_lpi_1_dfm_mx1);
  assign mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp = { _00836_, MulIn_data_sva_132[86:64] } * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4738" *) { _00837_, else_MulOp_data_2_lpi_1_dfm_2_30_0_1[22:0] };
  assign mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 = $signed(MulIn_data_sva_1[95:64]) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4747" *) $signed(else_MulOp_data_2_lpi_1_dfm_mx1);
  assign mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp = { _00839_, MulIn_data_sva_132[118:96] } * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4754" *) { _00840_, else_MulOp_data_3_lpi_1_dfm_2_30_0_1[22:0] };
  assign mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 = $signed(MulIn_data_sva_1[127:96]) * (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4763" *) $signed(else_MulOp_data_3_lpi_1_dfm_mx1);
  assign or_27_cse = cfg_precision != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4357" *) 2'b10;
  assign _00720_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4560" *) else_MulOp_data_0_lpi_1_dfm_mx0_30_0;
  assign _00721_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4561" *) else_MulOp_data_1_lpi_1_dfm_mx0_30_0;
  assign _00722_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4562" *) else_MulOp_data_2_lpi_1_dfm_mx0_30_0;
  assign _00723_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4563" *) else_MulOp_data_3_lpi_1_dfm_mx0_30_0;
  assign _00724_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4591" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva[63:31];
  assign _00725_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4619" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva[63:31];
  assign _00726_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4647" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva[63:31];
  assign _00727_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4675" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva[63:31];
  assign _00728_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4676" *) chn_mul_in_rsci_d_mxwt[30:0];
  assign _00729_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4677" *) chn_mul_in_rsci_d_mxwt[62:32];
  assign _00730_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4678" *) chn_mul_in_rsci_d_mxwt[94:64];
  assign _00731_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4679" *) chn_mul_in_rsci_d_mxwt[126:96];
  assign _00732_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4686" *) else_MulOp_data_0_lpi_1_dfm_mx0_30_0[22:0];
  assign _00733_ = else_MulOp_data_0_lpi_1_dfm_mx0_30_0[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4687" *) 8'b11111111;
  assign _00734_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4690" *) else_MulOp_data_1_lpi_1_dfm_mx0_30_0[22:0];
  assign _00735_ = else_MulOp_data_1_lpi_1_dfm_mx0_30_0[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4691" *) 8'b11111111;
  assign _00736_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4694" *) else_MulOp_data_2_lpi_1_dfm_mx0_30_0[22:0];
  assign _00737_ = else_MulOp_data_2_lpi_1_dfm_mx0_30_0[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4695" *) 8'b11111111;
  assign _00738_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4698" *) else_MulOp_data_3_lpi_1_dfm_mx0_30_0[22:0];
  assign _00739_ = else_MulOp_data_3_lpi_1_dfm_mx0_30_0[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4699" *) 8'b11111111;
  assign _00740_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4764" *) chn_mul_in_rsci_d_mxwt[22:0];
  assign _00741_ = chn_mul_in_rsci_d_mxwt[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4765" *) 8'b11111111;
  assign _00742_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4766" *) chn_mul_in_rsci_d_mxwt[54:32];
  assign _00743_ = chn_mul_in_rsci_d_mxwt[62:55] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4767" *) 8'b11111111;
  assign _00744_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4768" *) chn_mul_in_rsci_d_mxwt[86:64];
  assign _00745_ = chn_mul_in_rsci_d_mxwt[94:87] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4769" *) 8'b11111111;
  assign _00746_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4770" *) chn_mul_in_rsci_d_mxwt[118:96];
  assign _00747_ = chn_mul_in_rsci_d_mxwt[126:119] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4771" *) 8'b11111111;
  assign _00748_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4875" *) FpMul_8U_23U_o_expo_1_lpi_1_dfm;
  assign _00749_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4895" *) FpMul_8U_23U_o_expo_2_lpi_1_dfm;
  assign _00750_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4913" *) FpMul_8U_23U_o_expo_3_lpi_1_dfm;
  assign _00751_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4931" *) FpMul_8U_23U_o_expo_lpi_1_dfm;
  assign _00752_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4345" *) main_stage_v_3;
  assign _00753_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4345" *) _01024_;
  assign _00754_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4346" *) IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  assign _00755_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4347" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _00756_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4348" *) IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  assign _00757_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4350" *) IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  assign _00758_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4352" *) IsNaN_8U_23U_land_lpi_1_dfm_8;
  assign _00759_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4356" *) mux_7_itm;
  assign _00760_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4360" *) mux_12_itm;
  assign _00761_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4363" *) mux_17_itm;
  assign _00762_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4366" *) mux_22_itm;
  assign _00763_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4369" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _00764_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4371" *) and_dcpl_23;
  assign _00765_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4372" *) reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign _00766_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4373" *) main_stage_v_2;
  assign nor_319_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4373" *) _01026_;
  assign nor_320_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4375" *) _01028_;
  assign nor_315_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4379" *) _01030_;
  assign nor_316_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4381" *) _01032_;
  assign nor_311_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4385" *) _01034_;
  assign nor_312_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4387" *) _01036_;
  assign nor_307_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4391" *) _01038_;
  assign nor_308_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4393" *) _01040_;
  assign _00767_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4398" *) mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign nor_301_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4399" *) _01042_;
  assign nand_48_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4405" *) _00414_;
  assign nor_277_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4411" *) or_515_nl;
  assign _00768_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4412" *) mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign _00769_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4413" *) mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2;
  assign nor_282_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4413" *) _01045_;
  assign _00770_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4414" *) mux_tmp_48;
  assign _00771_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4417" *) mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign nor_264_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4418" *) _01046_;
  assign nor_348_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4419" *) _00846_;
  assign nor_267_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4420" *) _01047_;
  assign nand_45_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4424" *) _00416_;
  assign nor_241_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4430" *) or_523_nl;
  assign _00772_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4431" *) mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign _00773_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4432" *) mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2;
  assign nor_245_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4432" *) _01050_;
  assign _00774_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4433" *) mux_94_itm;
  assign _00775_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4436" *) mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign nor_227_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4437" *) _01051_;
  assign nor_347_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4438" *) _00848_;
  assign nor_230_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4439" *) _01052_;
  assign nand_42_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4443" *) _00417_;
  assign nor_204_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4449" *) or_531_nl;
  assign _00776_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4450" *) mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign _00777_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4451" *) mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2;
  assign nor_208_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4451" *) _01055_;
  assign _00778_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4452" *) mux_125_itm;
  assign _00779_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4455" *) mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign nor_190_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4456" *) _01057_;
  assign nor_346_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4457" *) _00850_;
  assign nor_193_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4458" *) _01058_;
  assign _00780_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4461" *) mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign nor_170_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4468" *) _01056_;
  assign _00781_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4470" *) mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2;
  assign nor_174_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4470" *) _01061_;
  assign _00782_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4471" *) mux_tmp_140;
  assign _00783_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4474" *) mux_tmp_46;
  assign _00784_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4475" *) and_20_tmp;
  assign _00785_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4475" *) _01062_;
  assign _00786_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4476" *) fsm_output[0];
  assign _00787_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4481" *) mux_160_nl;
  assign _00788_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4485" *) mux_168_nl;
  assign _00789_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4489" *) mux_173_nl;
  assign _00790_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4493" *) mux_178_nl;
  assign _00791_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4495" *) cfg_mul_bypass_rsci_d;
  assign nor_143_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4496" *) or_74_cse;
  assign _00792_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4497" *) or_dcpl_22;
  assign _00793_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4498" *) or_dcpl_27;
  assign _00794_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4500" *) _01064_;
  assign _00795_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4501" *) or_dcpl_37;
  assign _00796_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4502" *) or_dcpl_40;
  assign _00797_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4504" *) _01065_;
  assign _00798_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4505" *) or_dcpl_50;
  assign _00799_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4506" *) or_dcpl_53;
  assign _00800_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4508" *) _01066_;
  assign _00801_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4509" *) or_dcpl_63;
  assign _00802_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4510" *) or_dcpl_66;
  assign _00803_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4512" *) _01067_;
  assign _00804_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4513" *) IsNaN_8U_23U_land_1_lpi_1_dfm_4;
  assign _00806_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4517" *) IsNaN_8U_23U_land_2_lpi_1_dfm_4;
  assign _00808_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4521" *) IsNaN_8U_23U_land_3_lpi_1_dfm_4;
  assign _00810_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4525" *) IsNaN_8U_23U_land_lpi_1_dfm_4;
  assign nor_118_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4530" *) FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0;
  assign nor_117_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4534" *) FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0;
  assign nor_116_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4538" *) FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0;
  assign nor_115_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4542" *) _01071_;
  assign _00812_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4545" *) and_18_tmp;
  assign _00813_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4546" *) mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  assign _00814_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4548" *) mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  assign _00815_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4550" *) mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  assign _00816_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *) chn_mul_in_rsci_d_mxwt[31];
  assign _00817_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *) _01075_;
  assign _00818_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *) chn_mul_in_rsci_d_mxwt[63];
  assign _00819_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *) _01078_;
  assign _00820_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *) chn_mul_in_rsci_d_mxwt[95];
  assign _00821_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *) _01081_;
  assign _00822_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *) chn_mul_in_rsci_d_mxwt[127];
  assign _00823_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *) _01084_;
  assign IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4560" *) _00720_;
  assign IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4561" *) _00721_;
  assign IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4562" *) _00722_;
  assign IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4563" *) _00723_;
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4571" *) _00424_;
  assign _00824_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4589" *) FpMul_8U_23U_p_mant_p1_1_sva_mx1[47];
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4590" *) _00709_;
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4591" *) _00724_;
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4599" *) _00426_;
  assign _00825_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4617" *) FpMul_8U_23U_p_mant_p1_2_sva_mx1[47];
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4618" *) _00711_;
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4619" *) _00725_;
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4627" *) _00428_;
  assign _00826_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4645" *) FpMul_8U_23U_p_mant_p1_3_sva_mx1[47];
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4646" *) _00713_;
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4647" *) _00726_;
  assign FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4655" *) _00430_;
  assign _00827_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4673" *) FpMul_8U_23U_p_mant_p1_sva_mx1[47];
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4674" *) _00715_;
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4675" *) _00727_;
  assign IsZero_8U_23U_land_1_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4676" *) _00728_;
  assign IsZero_8U_23U_land_2_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4677" *) _00729_;
  assign IsZero_8U_23U_land_3_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4678" *) _00730_;
  assign IsZero_8U_23U_land_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4679" *) _00731_;
  assign _00828_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4680" *) cfg_mul_prelu_rsci_d;
  assign mul_mul_land_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4680" *) _01181_;
  assign mul_mul_land_3_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4681" *) _01182_;
  assign mul_mul_land_2_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4682" *) _01183_;
  assign mul_mul_land_1_lpi_1_dfm_mx1w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4683" *) _01184_;
  assign IsNaN_8U_23U_1_nor_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4686" *) _00732_;
  assign IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4687" *) _00805_;
  assign IsNaN_8U_23U_1_nor_1_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4690" *) _00734_;
  assign IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4691" *) _00807_;
  assign IsNaN_8U_23U_1_nor_2_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4694" *) _00736_;
  assign IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4695" *) _00809_;
  assign IsNaN_8U_23U_1_nor_3_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4698" *) _00738_;
  assign IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4699" *) _00811_;
  assign _00829_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4701" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  assign _00830_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4704" *) IsZero_8U_23U_land_1_lpi_1_dfm_6;
  assign _00831_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4705" *) IsZero_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _00832_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4717" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  assign _00833_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4720" *) IsZero_8U_23U_land_2_lpi_1_dfm_6;
  assign _00834_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4721" *) IsZero_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _00835_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4733" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  assign _00836_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4736" *) IsZero_8U_23U_land_3_lpi_1_dfm_6;
  assign _00837_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4737" *) IsZero_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _00838_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4749" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign _00839_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4752" *) IsZero_8U_23U_land_lpi_1_dfm_6;
  assign _00840_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4753" *) IsZero_8U_23U_1_land_lpi_1_dfm_6;
  assign _00841_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4764" *) _00740_;
  assign IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4765" *) _01186_;
  assign _00842_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4766" *) _00742_;
  assign IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4767" *) _01187_;
  assign _00843_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4768" *) _00744_;
  assign IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4769" *) _01188_;
  assign _00844_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4770" *) _00746_;
  assign IsNaN_8U_23U_land_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4771" *) _01189_;
  assign FpMul_8U_23U_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4779" *) _00012_;
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_4_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4781" *) _00013_;
  assign FpMul_8U_23U_FpMul_8U_23U_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4783" *) _01190_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_1_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4789" *) _01191_;
  assign mul_mul_else_unequal_tmp_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4792" *) and_dcpl_37;
  assign FpMul_8U_23U_nor_4_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4800" *) _00015_;
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_5_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4802" *) _00016_;
  assign FpMul_8U_23U_FpMul_8U_23U_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4804" *) _01192_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_2_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4810" *) _01193_;
  assign FpMul_8U_23U_nor_5_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4820" *) _00018_;
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_6_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4822" *) _00019_;
  assign FpMul_8U_23U_FpMul_8U_23U_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4824" *) _01194_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_3_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4830" *) _01195_;
  assign FpMul_8U_23U_nor_6_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4840" *) _00021_;
  assign FpMul_8U_23U_FpMul_8U_23U_FpMul_8U_23U_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4842" *) _00022_;
  assign FpMul_8U_23U_FpMul_8U_23U_nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4844" *) _01196_;
  assign IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_sva = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4850" *) _01197_;
  assign mul_mul_mul_mul_nor_6_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4853" *) _01198_;
  assign mul_mul_mul_mul_nor_4_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4854" *) _01199_;
  assign mul_mul_mul_mul_nor_2_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4855" *) _01200_;
  assign mul_mul_mul_mul_nor_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4856" *) _01201_;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4862" *) _00011_[22];
  assign FpMul_8U_23U_FpMul_8U_23U_nor_4_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4867" *) _01202_;
  assign _00845_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4875" *) _00748_;
  assign FpMul_8U_23U_is_inf_1_lpi_1_dfm_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4878" *) or_tmp_133;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4884" *) _00014_[22];
  assign _00847_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4895" *) _00749_;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4902" *) _00017_[22];
  assign _00849_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4913" *) _00750_;
  assign FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4920" *) _00020_[22];
  assign _00851_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4931" *) _00751_;
  assign _00852_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4980" *) _00447_;
  assign _00853_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4981" *) main_stage_v_1;
  assign _00854_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5498" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1086];
  assign _00855_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6014" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1086];
  assign _00856_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6530" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1086];
  assign _00857_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7046" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1086];
  assign _00858_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7088" *) mul_mul_land_lpi_1_dfm_6;
  assign _00859_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7091" *) mul_mul_land_1_lpi_1_dfm_6;
  assign _00860_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7094" *) mul_mul_land_3_lpi_1_dfm_6;
  assign _00861_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7097" *) mul_mul_land_2_lpi_1_dfm_6;
  assign _00862_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7112" *) mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7114" *) _05293_;
  assign nor_331_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7117" *) _05298_;
  assign _00863_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7127" *) mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign nor_326_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7129" *) _05306_;
  assign nor_327_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7132" *) _05311_;
  assign _00864_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7142" *) mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign nor_324_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7144" *) _05319_;
  assign nor_325_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7147" *) _05324_;
  assign _00865_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7156" *) mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign nor_321_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7157" *) _05334_;
  assign _00866_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7158" *) mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  assign nor_322_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7159" *) _05336_;
  assign nor_323_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7163" *) _05341_;
  assign nor_285_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7195" *) _05356_;
  assign nor_286_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7197" *) _05359_;
  assign nor_288_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7199" *) _05361_;
  assign nor_289_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7200" *) or_tmp_173;
  assign nor_283_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7207" *) _05365_;
  assign nor_284_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7209" *) _05368_;
  assign nor_248_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7222" *) _05378_;
  assign nor_249_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7224" *) _05381_;
  assign nor_251_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7226" *) _05383_;
  assign nor_252_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7228" *) _05384_;
  assign nor_246_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7234" *) _05388_;
  assign nor_247_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7236" *) _05391_;
  assign nor_211_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7250" *) _05401_;
  assign nor_212_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7252" *) _05404_;
  assign nor_214_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7254" *) _05406_;
  assign nor_215_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7256" *) _05407_;
  assign nor_209_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7262" *) _05411_;
  assign nor_210_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7264" *) _05414_;
  assign not_tmp_121 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7271" *) _00459_;
  assign nor_177_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7282" *) _05427_;
  assign nor_179_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7284" *) _05430_;
  assign nor_180_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7286" *) _05431_;
  assign nor_175_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7291" *) _05434_;
  assign nor_176_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7293" *) _05437_;
  assign _00867_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7296" *) _05441_;
  assign _00868_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7304" *) or_tmp_411;
  assign _00869_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7307" *) chn_mul_out_rsci_bawt;
  assign _00870_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7318" *) cfg_precision[0];
  assign _00871_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7319" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _00872_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7325" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _00873_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7329" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _00874_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7333" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _00875_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7342" *) cfg_precision[1];
  assign or_dcpl_96 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7359" *) _00463_;
  assign _00876_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7370" *) cfg_mul_src_rsci_d;
  assign _00877_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7387" *) _00469_;
  assign _00878_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7474" *) and_dcpl_26;
  assign _00879_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7482" *) chn_mul_op_rsci_ld_core_psct_mx0c1;
  assign _00880_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7490" *) main_stage_v_2_mx0c1;
  assign _00881_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7553" *) mux_9_nl;
  assign _00882_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7605" *) mux_14_nl;
  assign _00883_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7657" *) mux_19_nl;
  assign _00884_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7709" *) mux_24_nl;
  assign _00885_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7747" *) main_stage_v_3_mx0c1;
  assign _00886_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7866" *) mux_55_nl;
  assign _00887_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8003" *) mux_85_nl;
  assign _00888_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8140" *) mux_116_nl;
  assign _00889_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8267" *) mux_147_nl;
  assign _00890_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8277" *) mux_149_nl;
  assign _00891_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8383" *) main_stage_v_1_mx0c1;
  assign _00892_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8430" *) _05469_;
  assign _00893_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8439" *) or_tmp_461;
  assign _00894_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8539" *) _05471_;
  assign _00895_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8605" *) _05473_;
  assign _00896_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8670" *) _05475_;
  assign _00897_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8735" *) _05477_;
  assign _00898_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8768" *) and_dcpl_39;
  assign _00899_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8776" *) _05479_;
  assign _00900_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8804" *) _05483_;
  assign _00901_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8832" *) _05487_;
  assign _00902_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8860" *) _05491_;
  assign _00903_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8880" *) _05496_;
  assign _00904_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8902" *) _05498_;
  assign _00905_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8911" *) _05500_;
  assign _00906_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8932" *) _05503_;
  assign _00907_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8954" *) _05506_;
  assign _00908_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8975" *) or_dcpl_99;
  assign _00909_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8975" *) mux_164_nl;
  assign _00910_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8983" *) _05508_;
  assign _00911_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8991" *) or_dcpl_102;
  assign _00912_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8991" *) mux_172_nl;
  assign _00913_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8999" *) _05509_;
  assign _00914_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9007" *) or_dcpl_105;
  assign _00915_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9007" *) mux_177_nl;
  assign _00916_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9015" *) _05510_;
  assign _00917_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9023" *) or_dcpl_108;
  assign _00918_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9023" *) mux_182_nl;
  assign _00919_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9031" *) _05511_;
  assign _00920_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9079" *) _05512_;
  assign _00921_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *) _05517_;
  assign _00922_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9098" *) _05520_;
  assign _00923_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *) _05525_;
  assign _00924_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9117" *) _05528_;
  assign _00925_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *) _05533_;
  assign _00926_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9136" *) _05536_;
  assign _00927_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9146" *) _05541_;
  assign _00928_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9155" *) _05544_;
  assign _00929_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9161" *) _05545_;
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9161" *) _05546_;
  assign _00930_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9169" *) _05547_;
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9169" *) _05548_;
  assign _00931_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9176" *) _05549_;
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9176" *) _05550_;
  assign _00932_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9184" *) _05551_;
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9184" *) _05552_;
  assign _00933_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9191" *) _05553_;
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9191" *) _05554_;
  assign _00934_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9199" *) _05555_;
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9199" *) _05556_;
  assign _00935_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9205" *) _05557_;
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9206" *) _05558_;
  assign _00936_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9213" *) _05559_;
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9214" *) _05560_;
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9220" *) _00003_;
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9223" *) _00004_;
  assign nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9224" *) _05561_;
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9229" *) _00023_;
  assign mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9232" *) _00024_;
  assign _00937_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9233" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9238" *) _00005_;
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9241" *) _00006_;
  assign nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9242" *) _05562_;
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9247" *) _00025_;
  assign mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9250" *) _00026_;
  assign _00938_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9251" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9256" *) _00007_;
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9259" *) _00008_;
  assign nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9260" *) _05563_;
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9265" *) _00027_;
  assign mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9268" *) _00028_;
  assign _00939_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9269" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9274" *) _00009_;
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9277" *) _00010_;
  assign nor_6_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9278" *) _05564_;
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9283" *) _00029_;
  assign mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9286" *) _00030_;
  assign _00940_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9287" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign nor_299_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9320" *) _05585_;
  assign _00941_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9323" *) FpMul_8U_23U_lor_6_lpi_1_dfm_6;
  assign _00942_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9327" *) or_tmp_128;
  assign _00943_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9331" *) _05592_;
  assign nor_300_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9335" *) _05593_;
  assign _00944_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9338" *) _05362_;
  assign _00945_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9340" *) or_tmp_132;
  assign nor_304_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9340" *) _05594_;
  assign _00946_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9343" *) _00618_;
  assign nor_303_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9347" *) _05595_;
  assign nor_296_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9350" *) _05599_;
  assign _00947_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9351" *) mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign nor_297_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9353" *) _05603_;
  assign _00948_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9357" *) _00619_;
  assign nor_298_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9357" *) _05606_;
  assign nor_292_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9371" *) _05613_;
  assign _00949_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9375" *) _00620_;
  assign nor_294_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9375" *) _05616_;
  assign nor_290_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9378" *) _05617_;
  assign _00950_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9380" *) mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign nor_291_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9380" *) _05618_;
  assign nor_276_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9388" *) _05624_;
  assign nor_278_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9390" *) _05626_;
  assign nand_15_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9393" *) _00621_;
  assign _00951_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9394" *) FpMul_8U_23U_FpMul_8U_23U_and_itm;
  assign nor_275_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9400" *) _05628_;
  assign _00952_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *) FpMul_8U_23U_FpMul_8U_23U_and_itm_2;
  assign _00953_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *) _05630_;
  assign _00954_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *) _05631_;
  assign nor_279_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *) _05632_;
  assign nor_269_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9407" *) _05639_;
  assign nor_271_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9410" *) _05646_;
  assign nor_272_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9416" *) _05653_;
  assign nor_273_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9420" *) _05661_;
  assign _00955_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9426" *) FpMul_8U_23U_lor_7_lpi_1_dfm_6;
  assign _00956_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9431" *) or_tmp_216;
  assign _00957_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9435" *) _05672_;
  assign nor_263_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9440" *) _05673_;
  assign _00958_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9441" *) mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign nor_268_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9441" *) _05674_;
  assign _00959_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9444" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_4;
  assign nand_20_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9447" *) _00625_;
  assign nor_266_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9451" *) _05676_;
  assign nor_260_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9454" *) _05680_;
  assign _00960_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9455" *) mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign nor_261_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9457" *) _05684_;
  assign _00961_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9461" *) _00626_;
  assign nor_262_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9461" *) _05687_;
  assign nor_255_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9475" *) _05694_;
  assign _00962_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9476" *) _05675_;
  assign nor_257_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9479" *) _05702_;
  assign nor_253_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9482" *) _05703_;
  assign nor_254_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9484" *) _05704_;
  assign nor_238_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9490" *) _05706_;
  assign nor_240_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9492" *) _05709_;
  assign nor_242_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9494" *) _05712_;
  assign nand_22_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9497" *) _00627_;
  assign _00963_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9498" *) FpMul_8U_23U_FpMul_8U_23U_and_12_itm;
  assign nor_239_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9501" *) _05715_;
  assign _00964_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9504" *) _05385_;
  assign _00965_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9507" *) FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2;
  assign _00966_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9507" *) _05717_;
  assign _00967_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9508" *) _05718_;
  assign nor_243_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9508" *) _05719_;
  assign nor_232_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9512" *) _05725_;
  assign nor_234_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9515" *) _05731_;
  assign nor_235_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9521" *) _05737_;
  assign nor_236_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9525" *) _05745_;
  assign _00968_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9531" *) FpMul_8U_23U_lor_8_lpi_1_dfm_6;
  assign _00969_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9536" *) or_tmp_296;
  assign _00970_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9540" *) _05756_;
  assign nor_226_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9545" *) _05757_;
  assign _00971_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9546" *) mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign nor_231_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9546" *) _05758_;
  assign _00972_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9549" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_4;
  assign nand_27_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9552" *) _00631_;
  assign nor_229_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9556" *) _05760_;
  assign nor_223_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9559" *) _05764_;
  assign _00973_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9560" *) mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign nor_224_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9562" *) _05768_;
  assign _00974_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9566" *) _00632_;
  assign nor_225_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9566" *) _05771_;
  assign nor_218_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9580" *) _05778_;
  assign _00975_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9581" *) _05759_;
  assign nor_220_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9584" *) _05786_;
  assign nor_216_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9587" *) _05787_;
  assign nor_217_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9589" *) _05788_;
  assign nor_201_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9595" *) _05790_;
  assign nor_203_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9597" *) _05793_;
  assign nor_205_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9599" *) _05796_;
  assign nand_29_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9602" *) _00633_;
  assign _00976_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9603" *) FpMul_8U_23U_FpMul_8U_23U_and_13_itm;
  assign nor_202_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9606" *) _05799_;
  assign _00977_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9609" *) _05408_;
  assign _00978_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9612" *) FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2;
  assign _00979_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9612" *) _05801_;
  assign _00980_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9613" *) _05802_;
  assign nor_206_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9613" *) _05803_;
  assign nor_195_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9617" *) _05809_;
  assign nor_197_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9620" *) _05815_;
  assign nor_198_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9626" *) _05821_;
  assign nor_199_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9630" *) _05829_;
  assign _00981_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9636" *) FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  assign _00982_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9641" *) or_tmp_376;
  assign _00983_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9645" *) _05840_;
  assign nor_189_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9650" *) _05841_;
  assign _00984_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9651" *) mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign nor_194_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9651" *) or_424_nl;
  assign _00985_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9654" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_4;
  assign nand_34_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9657" *) _00637_;
  assign nor_192_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9661" *) _05843_;
  assign nor_186_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9664" *) _05847_;
  assign _00986_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9665" *) mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign nor_187_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9667" *) _05851_;
  assign _00987_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9671" *) _00638_;
  assign nor_188_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9671" *) _05854_;
  assign nor_181_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9685" *) _05861_;
  assign _00988_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9686" *) _05842_;
  assign nor_183_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9689" *) _05869_;
  assign nor_167_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9701" *) _05871_;
  assign nor_169_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9703" *) _05874_;
  assign nor_171_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9705" *) _05877_;
  assign nand_36_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9708" *) _00639_;
  assign _00989_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9709" *) FpMul_8U_23U_FpMul_8U_23U_and_14_itm;
  assign nor_168_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9712" *) _05880_;
  assign _00990_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9715" *) or_435_nl;
  assign _00991_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9718" *) FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2;
  assign _00992_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9718" *) _05882_;
  assign _00993_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9719" *) _05883_;
  assign nor_172_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9719" *) _05884_;
  assign nor_161_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9723" *) _05890_;
  assign nor_163_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9726" *) _05896_;
  assign nor_164_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9732" *) _05902_;
  assign nor_165_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9736" *) _05910_;
  assign nor_144_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9741" *) _05913_;
  assign _00000_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9748" *) FpMul_8U_23U_p_mant_p1_1_sva[47];
  assign nor_142_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9761" *) _05923_;
  assign _00001_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9766" *) FpMul_8U_23U_p_mant_p1_2_sva[47];
  assign nor_140_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9779" *) _05930_;
  assign _00002_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9784" *) FpMul_8U_23U_p_mant_p1_3_sva[47];
  assign nor_342_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9797" *) _05935_;
  assign _00994_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9801" *) mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign nor_136_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9812" *) _05938_;
  assign nor_137_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9815" *) _05942_;
  assign nor_138_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9820" *) _05947_;
  assign nor_134_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9823" *) _05948_;
  assign nor_135_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9825" *) _05951_;
  assign nor_131_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9830" *) _05953_;
  assign nor_132_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9833" *) _05957_;
  assign nor_133_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9838" *) _05962_;
  assign nor_129_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9841" *) _05963_;
  assign nor_130_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9843" *) _05966_;
  assign nor_126_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9848" *) _05968_;
  assign nor_127_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9851" *) _05972_;
  assign nor_128_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9856" *) _05977_;
  assign nor_124_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9859" *) _05978_;
  assign nor_125_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9861" *) _05981_;
  assign nor_121_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9866" *) _05983_;
  assign nor_122_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9869" *) _05987_;
  assign nor_123_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9874" *) _05992_;
  assign nor_119_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9877" *) _05993_;
  assign nor_120_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9879" *) _05996_;
  assign nor_159_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9881" *) _05997_;
  assign _00995_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9883" *) or_tmp_1;
  assign nor_157_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9890" *) _06002_;
  assign _00996_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9892" *) or_tmp_15;
  assign nor_155_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9899" *) _06007_;
  assign _00997_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9901" *) or_tmp_29;
  assign nor_153_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9910" *) _06012_;
  assign _00998_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9912" *) or_tmp_46;
  assign _00999_ = _00374_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) _00382_;
  assign _01000_ = _00375_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) _00383_;
  assign _01001_ = _00376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) _00384_;
  assign _01002_ = _00377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) _00385_;
  assign _01003_ = _00378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) _00386_;
  assign _01004_ = _00379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) _00387_;
  assign _01005_ = _00380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) _00388_;
  assign _01006_ = _00381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10004" *) _00389_;
  assign _01007_ = _00999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) _00390_;
  assign _01008_ = _01000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) _00391_;
  assign _01009_ = _01001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) _00392_;
  assign _01010_ = _01002_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) _00393_;
  assign _01011_ = _01003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) _00394_;
  assign _01012_ = _01004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) _00395_;
  assign _01013_ = _01005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) _00396_;
  assign _01014_ = _01006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10005" *) _00397_;
  assign _01015_ = _01007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) _00398_;
  assign _01016_ = _01008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) _00399_;
  assign _01017_ = _01009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) _00400_;
  assign _01018_ = _01010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) _00401_;
  assign _01019_ = _01011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) _00402_;
  assign _01020_ = _01012_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) _00403_;
  assign _01021_ = _01013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) _00404_;
  assign _01022_ = _01014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10006" *) _00405_;
  assign _01023_ = _00407_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4344" *) and_dcpl_22;
  assign _01024_ = and_dcpl_23 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4345" *) _00752_;
  assign IsZero_8U_23U_1_aelse_IsZero_8U_23U_1_aelse_or_3_cse = and_dcpl_38 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4355" *) and_dcpl_39;
  assign or_74_cse = _00765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4372" *) chn_mul_out_rsci_bawt;
  assign _01025_ = _00766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4373" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _01026_ = _01025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4373" *) or_tmp_59;
  assign or_tmp_173 = _00752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4374" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _01027_ = or_tmp_173 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4375" *) mul_mul_land_1_lpi_1_dfm_6;
  assign _01028_ = _01027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4375" *) mul_mul_land_1_lpi_1_dfm_st_5;
  assign _01029_ = _00766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4379" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _01030_ = _01029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4379" *) or_tmp_75;
  assign _01031_ = or_tmp_173 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4381" *) mul_mul_land_2_lpi_1_dfm_6;
  assign _01032_ = _01031_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4381" *) mul_mul_land_2_lpi_1_dfm_st_5;
  assign _01033_ = _00766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4385" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _01034_ = _01033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4385" *) or_tmp_91;
  assign _01035_ = or_tmp_173 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4387" *) mul_mul_land_3_lpi_1_dfm_6;
  assign _01036_ = _01035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4387" *) mul_mul_land_3_lpi_1_dfm_st_5;
  assign _01037_ = _00766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4391" *) mul_mul_land_lpi_1_dfm_5;
  assign _01038_ = _01037_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4391" *) or_tmp_107;
  assign _01039_ = or_tmp_173 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4393" *) mul_mul_land_lpi_1_dfm_6;
  assign _01040_ = _01039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4393" *) mul_mul_land_lpi_1_dfm_st_5;
  assign _01041_ = FpMul_8U_23U_lor_6_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4399" *) _00767_;
  assign _01042_ = _01041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4399" *) mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign _01043_ = and_dcpl_46 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4401" *) and_dcpl_48;
  assign _01044_ = _01043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4401" *) and_dcpl_50;
  assign FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_3_cse = _01044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4401" *) and_dcpl_51;
  assign FpMul_8U_23U_else_2_else_if_FpMul_8U_23U_else_2_else_if_or_7_cse = and_dcpl_52 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4403" *) and_dcpl_47;
  assign or_515_nl = _00767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4411" *) mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign or_743_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4412" *) _00768_;
  assign _01045_ = _00769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4413" *) mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2;
  assign or_523_nl = _00771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4418" *) mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign _01046_ = or_523_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4418" *) FpMul_8U_23U_lor_7_lpi_1_dfm_6;
  assign _00846_ = FpMul_8U_23U_lor_7_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4419" *) FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2;
  assign _01047_ = nor_348_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4420" *) mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2;
  assign _01048_ = and_dcpl_54 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4422" *) and_dcpl_55;
  assign _01049_ = _01048_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4422" *) and_dcpl_57;
  assign FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_2_cse = _01049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4422" *) and_dcpl_58;
  assign or_744_nl = FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4431" *) _00772_;
  assign _01050_ = _00773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4432" *) mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2;
  assign or_531_nl = _00775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4437" *) mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign _01051_ = or_531_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4437" *) FpMul_8U_23U_lor_8_lpi_1_dfm_6;
  assign _00848_ = FpMul_8U_23U_lor_8_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4438" *) FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2;
  assign _01052_ = nor_347_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4439" *) mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2;
  assign _01053_ = and_dcpl_60 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4441" *) and_dcpl_61;
  assign _01054_ = _01053_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4441" *) and_dcpl_63;
  assign FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_1_cse = _01054_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4441" *) and_dcpl_64;
  assign or_745_nl = FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4450" *) _00776_;
  assign _01055_ = _00777_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4451" *) mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2;
  assign _01056_ = _00779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4456" *) mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign _01057_ = _01056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4456" *) FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  assign _00850_ = FpMul_8U_23U_lor_1_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4457" *) FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2;
  assign _01058_ = nor_346_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4458" *) mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2;
  assign _01059_ = and_dcpl_66 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4460" *) and_dcpl_67;
  assign _01060_ = _01059_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4460" *) and_dcpl_69;
  assign FpMul_8U_23U_p_expo_FpMul_8U_23U_p_expo_or_cse = _01060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4460" *) and_dcpl_70;
  assign or_430_cse = _00780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4462" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign _01061_ = _00781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4470" *) mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2;
  assign _01062_ = _00784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4475" *) fsm_output[0];
  assign IsNaN_8U_23U_aelse_IsNaN_8U_23U_aelse_or_3_cse = and_dcpl_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4477" *) and_dcpl_6;
  assign or_467_nl = mul_mul_land_1_lpi_1_dfm_mx1w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4478" *) cfg_mul_bypass_rsci_d;
  assign or_480_nl = mul_mul_land_2_lpi_1_dfm_mx1w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4482" *) cfg_mul_bypass_rsci_d;
  assign or_488_nl = mul_mul_land_3_lpi_1_dfm_mx1w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4486" *) cfg_mul_bypass_rsci_d;
  assign or_496_nl = mul_mul_land_lpi_1_dfm_mx1w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4490" *) cfg_mul_bypass_rsci_d;
  assign _01063_ = or_dcpl_26 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4500" *) and_dcpl_37;
  assign _01064_ = _01063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4500" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign _01065_ = _01063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4504" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign _01066_ = _01063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4508" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign _01067_ = _01063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4512" *) mul_mul_land_lpi_1_dfm_st_4;
  assign or_dcpl_75 = IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4530" *) mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0 = or_dcpl_75 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4530" *) IsZero_8U_23U_land_1_lpi_1_dfm_4;
  assign _01068_ = FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4531" *) or_27_cse;
  assign or_dcpl_81 = IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4534" *) mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0 = or_dcpl_81 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4534" *) IsZero_8U_23U_land_2_lpi_1_dfm_4;
  assign _01069_ = FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4535" *) or_27_cse;
  assign or_dcpl_87 = IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4538" *) mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0 = or_dcpl_87 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4538" *) IsZero_8U_23U_land_3_lpi_1_dfm_4;
  assign _01070_ = FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4539" *) or_27_cse;
  assign or_dcpl_93 = IsZero_8U_23U_land_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4542" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp;
  assign _01071_ = or_dcpl_93 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4542" *) mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign _01072_ = _01071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4544" *) or_27_cse;
  assign or_468_cse = _00812_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4545" *) or_27_cse;
  assign or_469_cse = _00813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4547" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st;
  assign or_482_cse = _00814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4549" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st;
  assign or_490_cse = _00815_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4551" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st;
  assign _01073_ = _00420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *) cfg_mul_bypass_rsci_d;
  assign _01074_ = _01073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *) or_dcpl_110;
  assign _01075_ = _01074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4553" *) fsm_output[0];
  assign _01076_ = _00421_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *) cfg_mul_bypass_rsci_d;
  assign _01077_ = _01076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *) or_dcpl_110;
  assign _01078_ = _01077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4555" *) fsm_output[0];
  assign _01079_ = _00422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *) cfg_mul_bypass_rsci_d;
  assign _01080_ = _01079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *) or_dcpl_110;
  assign _01081_ = _01080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4557" *) fsm_output[0];
  assign _01082_ = _00423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *) cfg_mul_bypass_rsci_d;
  assign _01083_ = _01082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *) or_dcpl_110;
  assign _01084_ = _01083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4559" *) fsm_output[0];
  assign _01085_ = _00425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4576" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[0];
  assign _01086_ = _01085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4577" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[1];
  assign _01087_ = _01086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4577" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[2];
  assign _01088_ = _01087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4578" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[3];
  assign _01089_ = _01088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4578" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[4];
  assign _01090_ = _01089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4579" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[5];
  assign _01091_ = _01090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4579" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[6];
  assign _01092_ = _01091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4580" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[7];
  assign _01093_ = _01092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4580" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[8];
  assign _01094_ = _01093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4581" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[9];
  assign _01095_ = _01094_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4581" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[10];
  assign _01096_ = _01095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4582" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[11];
  assign _01097_ = _01096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4582" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[12];
  assign _01098_ = _01097_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4583" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[13];
  assign _01099_ = _01098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4583" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[14];
  assign _01100_ = _01099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4584" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[15];
  assign _01101_ = _01100_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4584" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[16];
  assign _01102_ = _01101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4585" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[17];
  assign _01103_ = _01102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4585" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[18];
  assign _01104_ = _01103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4586" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[19];
  assign _01105_ = _01104_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4586" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[20];
  assign _01106_ = _01105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4587" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[21];
  assign _01107_ = _01106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4587" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[23];
  assign _01108_ = mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4589" *) _00824_;
  assign _01109_ = _00427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4604" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[0];
  assign _01110_ = _01109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4605" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[1];
  assign _01111_ = _01110_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4605" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[2];
  assign _01112_ = _01111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4606" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[3];
  assign _01113_ = _01112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4606" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[4];
  assign _01114_ = _01113_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4607" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[5];
  assign _01115_ = _01114_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4607" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[6];
  assign _01116_ = _01115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4608" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[7];
  assign _01117_ = _01116_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4608" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[8];
  assign _01118_ = _01117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4609" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[9];
  assign _01119_ = _01118_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4609" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[10];
  assign _01120_ = _01119_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4610" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[11];
  assign _01121_ = _01120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4610" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[12];
  assign _01122_ = _01121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4611" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[13];
  assign _01123_ = _01122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4611" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[14];
  assign _01124_ = _01123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4612" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[15];
  assign _01125_ = _01124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4612" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[16];
  assign _01126_ = _01125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4613" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[17];
  assign _01127_ = _01126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4613" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[18];
  assign _01128_ = _01127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4614" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[19];
  assign _01129_ = _01128_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4614" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[20];
  assign _01130_ = _01129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4615" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[21];
  assign _01131_ = _01130_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4615" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[23];
  assign _01132_ = mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4617" *) _00825_;
  assign _01133_ = _00429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4632" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[0];
  assign _01134_ = _01133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4633" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[1];
  assign _01135_ = _01134_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4633" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[2];
  assign _01136_ = _01135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4634" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[3];
  assign _01137_ = _01136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4634" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[4];
  assign _01138_ = _01137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4635" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[5];
  assign _01139_ = _01138_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4635" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[6];
  assign _01140_ = _01139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4636" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[7];
  assign _01141_ = _01140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4636" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[8];
  assign _01142_ = _01141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4637" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[9];
  assign _01143_ = _01142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4637" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[10];
  assign _01144_ = _01143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4638" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[11];
  assign _01145_ = _01144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4638" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[12];
  assign _01146_ = _01145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4639" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[13];
  assign _01147_ = _01146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4639" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[14];
  assign _01148_ = _01147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4640" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[15];
  assign _01149_ = _01148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4640" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[16];
  assign _01150_ = _01149_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4641" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[17];
  assign _01151_ = _01150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4641" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[18];
  assign _01152_ = _01151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4642" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[19];
  assign _01153_ = _01152_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4642" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[20];
  assign _01154_ = _01153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4643" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[21];
  assign _01155_ = _01154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4643" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[23];
  assign _01156_ = mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4645" *) _00826_;
  assign _01157_ = _00431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4660" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[0];
  assign _01158_ = _01157_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4661" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[1];
  assign _01159_ = _01158_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4661" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[2];
  assign _01160_ = _01159_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4662" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[3];
  assign _01161_ = _01160_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4662" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[4];
  assign _01162_ = _01161_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4663" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[5];
  assign _01163_ = _01162_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4663" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[6];
  assign _01164_ = _01163_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4664" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[7];
  assign _01165_ = _01164_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4664" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[8];
  assign _01166_ = _01165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4665" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[9];
  assign _01167_ = _01166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4665" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[10];
  assign _01168_ = _01167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4666" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[11];
  assign _01169_ = _01168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4666" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[12];
  assign _01170_ = _01169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4667" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[13];
  assign _01171_ = _01170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4667" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[14];
  assign _01172_ = _01171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4668" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[15];
  assign _01173_ = _01172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4668" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[16];
  assign _01174_ = _01173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4669" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[17];
  assign _01175_ = _01174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4669" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[18];
  assign _01176_ = _01175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4670" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[19];
  assign _01177_ = _01176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4670" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[20];
  assign _01178_ = _01177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4671" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[21];
  assign _01179_ = _01178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4671" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[23];
  assign _01180_ = mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4673" *) _00827_;
  assign _01181_ = chn_mul_in_rsci_d_mxwt[127] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4680" *) _00828_;
  assign _01182_ = chn_mul_in_rsci_d_mxwt[95] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4681" *) _00828_;
  assign _01183_ = chn_mul_in_rsci_d_mxwt[63] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4682" *) _00828_;
  assign _01184_ = chn_mul_in_rsci_d_mxwt[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4683" *) _00828_;
  assign _00805_ = IsNaN_8U_23U_1_nor_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4687" *) _00733_;
  assign _00807_ = IsNaN_8U_23U_1_nor_1_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4691" *) _00735_;
  assign _00809_ = IsNaN_8U_23U_1_nor_2_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4695" *) _00737_;
  assign _01185_ = mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl[9] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4697" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp;
  assign FpMul_8U_23U_lor_1_lpi_1_dfm_mx0w0 = _01185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4697" *) IsZero_8U_23U_land_lpi_1_dfm_4;
  assign _00811_ = IsNaN_8U_23U_1_nor_3_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4699" *) _00739_;
  assign _01186_ = _00841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4765" *) _00741_;
  assign _01187_ = _00842_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4767" *) _00743_;
  assign _01188_ = _00843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4769" *) _00745_;
  assign _01189_ = _00844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4771" *) _00747_;
  assign or_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4775" *) _00769_;
  assign _01190_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4783" *) IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  assign _01191_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_64_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4789" *) mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  assign or_840_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4796" *) _00773_;
  assign _01192_ = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4804" *) IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  assign _01193_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_64_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4810" *) mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  assign or_841_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4816" *) _00777_;
  assign _01194_ = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4824" *) IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  assign _01195_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_64_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4830" *) mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  assign or_842_nl = FpMantWidthDec_8U_47U_23U_0U_0U_if_1_unequal_tmp_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4836" *) _00781_;
  assign _01196_ = IsNaN_8U_23U_1_land_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4844" *) IsNaN_8U_23U_land_lpi_1_dfm_8;
  assign _01197_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_64_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4850" *) mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  assign _01198_ = mul_mul_else_unequal_tmp_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4853" *) mul_mul_land_lpi_1_dfm_6;
  assign _01199_ = mul_mul_else_unequal_tmp_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4854" *) mul_mul_land_3_lpi_1_dfm_6;
  assign _01200_ = mul_mul_else_unequal_tmp_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4855" *) mul_mul_land_2_lpi_1_dfm_6;
  assign _01201_ = mul_mul_else_unequal_tmp_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4856" *) mul_mul_land_1_lpi_1_dfm_6;
  assign _01202_ = mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4867" *) FpMul_8U_23U_is_inf_1_lpi_1_dfm_2;
  assign FpMul_8U_23U_or_4_nl = _00432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4869" *) FpMul_8U_23U_is_inf_1_lpi_1_dfm_2;
  assign FpMul_8U_23U_lor_9_lpi_1_dfm = _00845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4876" *) FpMul_8U_23U_lor_6_lpi_1_dfm_7;
  assign or_tmp_133 = FpMul_8U_23U_FpMul_8U_23U_and_itm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4878" *) FpMul_8U_23U_lor_6_lpi_1_dfm_7;
  assign FpMul_8U_23U_or_5_nl = _00434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4889" *) nor_348_cse;
  assign FpMul_8U_23U_lor_10_lpi_1_dfm = _00847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4896" *) FpMul_8U_23U_lor_7_lpi_1_dfm_7;
  assign FpMul_8U_23U_or_6_nl = _00436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4907" *) nor_347_cse;
  assign FpMul_8U_23U_lor_11_lpi_1_dfm = _00849_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4914" *) FpMul_8U_23U_lor_8_lpi_1_dfm_7;
  assign FpMul_8U_23U_or_7_nl = _00438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4925" *) nor_346_cse;
  assign FpMul_8U_23U_lor_2_lpi_1_dfm = _00851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4932" *) FpMul_8U_23U_lor_1_lpi_1_dfm_7;
  assign or_11_cse = chn_mul_op_rsci_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4980" *) _00852_;
  assign or_12_cse = cfg_truncate_rsc_triosy_obj_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4981" *) _00853_;
  assign or_13_cse = cfg_mul_op_rsc_triosy_obj_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4982" *) _00853_;
  assign or_14_cse = cfg_mul_src_rsc_triosy_obj_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4983" *) _00853_;
  assign or_15_cse = cfg_mul_prelu_rsc_triosy_obj_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4984" *) _00853_;
  assign or_16_cse = cfg_mul_bypass_rsc_triosy_obj_bawt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4985" *) _00853_;
  assign _01203_ = IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4988" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1];
  assign _01204_ = _01203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4988" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[2];
  assign _01205_ = _01204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4989" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[3];
  assign _01206_ = _01205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4989" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[4];
  assign _01207_ = _01206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4990" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[5];
  assign _01208_ = _01207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4990" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[6];
  assign _01209_ = _01208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4991" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[7];
  assign _01210_ = _01209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4991" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[8];
  assign _01211_ = _01210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4992" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[9];
  assign _01212_ = _01211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4992" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[10];
  assign _01213_ = _01212_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4993" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[11];
  assign _01214_ = _01213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4993" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[12];
  assign _01215_ = _01214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4994" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[13];
  assign _01216_ = _01215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4994" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[14];
  assign _01217_ = _01216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4995" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[15];
  assign _01218_ = _01217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4995" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[16];
  assign _01219_ = _01218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4996" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[17];
  assign _01220_ = _01219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4996" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[18];
  assign _01221_ = _01220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4997" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[19];
  assign _01222_ = _01221_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4997" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[20];
  assign _01223_ = _01222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4998" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[21];
  assign _01224_ = _01223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4998" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[22];
  assign _01225_ = _01224_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4999" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[23];
  assign _01226_ = _01225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4999" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[24];
  assign _01227_ = _01226_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5000" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[25];
  assign _01228_ = _01227_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5000" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[26];
  assign _01229_ = _01228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5001" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[27];
  assign _01230_ = _01229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5001" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[28];
  assign _01231_ = _01230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5002" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[29];
  assign _01232_ = _01231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5002" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[30];
  assign _01233_ = _01232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5003" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[31];
  assign _01234_ = _01233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5003" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[32];
  assign _01235_ = _01234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5004" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[33];
  assign _01236_ = _01235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5004" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[34];
  assign _01237_ = _01236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5005" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[35];
  assign _01238_ = _01237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5005" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[36];
  assign _01239_ = _01238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5006" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[37];
  assign _01240_ = _01239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5006" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[38];
  assign _01241_ = _01240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5007" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[39];
  assign _01242_ = _01241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5007" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[40];
  assign _01243_ = _01242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5008" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[41];
  assign _01244_ = _01243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5008" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[42];
  assign _01245_ = _01244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5009" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[43];
  assign _01246_ = _01245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5009" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[44];
  assign _01247_ = _01246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5010" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[45];
  assign _01248_ = _01247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5010" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[46];
  assign _01249_ = _01248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5011" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[47];
  assign _01250_ = _01249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5011" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[48];
  assign _01251_ = _01250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5012" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[49];
  assign _01252_ = _01251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5012" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[50];
  assign _01253_ = _01252_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5013" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[51];
  assign _01254_ = _01253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5013" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[52];
  assign _01255_ = _01254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5014" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[53];
  assign _01256_ = _01255_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5014" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[54];
  assign _01257_ = _01256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5015" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[55];
  assign _01258_ = _01257_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5015" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[56];
  assign _01259_ = _01258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5016" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[57];
  assign _01260_ = _01259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5016" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[58];
  assign _01261_ = _01260_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5017" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[59];
  assign _01262_ = _01261_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5017" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[60];
  assign _01263_ = _01262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5018" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[61];
  assign _01264_ = _01263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5018" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[62];
  assign _01265_ = _01264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5019" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[63];
  assign _01266_ = _01265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5019" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[64];
  assign _01267_ = _01266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5020" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[65];
  assign _01268_ = _01267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5020" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[66];
  assign _01269_ = _01268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5021" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[67];
  assign _01270_ = _01269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5021" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[68];
  assign _01271_ = _01270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5022" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[69];
  assign _01272_ = _01271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5022" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[70];
  assign _01273_ = _01272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5023" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[71];
  assign _01274_ = _01273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5023" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[72];
  assign _01275_ = _01274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5024" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[73];
  assign _01276_ = _01275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5024" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[74];
  assign _01277_ = _01276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5025" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[75];
  assign _01278_ = _01277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5025" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[76];
  assign _01279_ = _01278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5026" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[77];
  assign _01280_ = _01279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5026" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[78];
  assign _01281_ = _01280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5027" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[79];
  assign _01282_ = _01281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5027" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[80];
  assign _01283_ = _01282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5028" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[81];
  assign _01284_ = _01283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5028" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[82];
  assign _01285_ = _01284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5029" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[83];
  assign _01286_ = _01285_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5029" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[84];
  assign _01287_ = _01286_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5030" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[85];
  assign _01288_ = _01287_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5030" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[86];
  assign _01289_ = _01288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5031" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[87];
  assign _01290_ = _01289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5031" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[88];
  assign _01291_ = _01290_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5032" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[89];
  assign _01292_ = _01291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5032" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[90];
  assign _01293_ = _01292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5033" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[91];
  assign _01294_ = _01293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5033" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[92];
  assign _01295_ = _01294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5034" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[93];
  assign _01296_ = _01295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5034" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[94];
  assign _01297_ = _01296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5035" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[95];
  assign _01298_ = _01297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5035" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[96];
  assign _01299_ = _01298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5036" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[97];
  assign _01300_ = _01299_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5036" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[98];
  assign _01301_ = _01300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5037" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[99];
  assign _01302_ = _01301_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5037" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[100];
  assign _01303_ = _01302_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5038" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[101];
  assign _01304_ = _01303_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5038" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[102];
  assign _01305_ = _01304_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5039" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[103];
  assign _01306_ = _01305_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5039" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[104];
  assign _01307_ = _01306_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5040" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[105];
  assign _01308_ = _01307_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5040" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[106];
  assign _01309_ = _01308_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5041" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[107];
  assign _01310_ = _01309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5041" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[108];
  assign _01311_ = _01310_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5042" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[109];
  assign _01312_ = _01311_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5042" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[110];
  assign _01313_ = _01312_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5043" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[111];
  assign _01314_ = _01313_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5043" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[112];
  assign _01315_ = _01314_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5044" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[113];
  assign _01316_ = _01315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5044" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[114];
  assign _01317_ = _01316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5045" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[115];
  assign _01318_ = _01317_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5045" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[116];
  assign _01319_ = _01318_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5046" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[117];
  assign _01320_ = _01319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5046" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[118];
  assign _01321_ = _01320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5047" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[119];
  assign _01322_ = _01321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5047" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[120];
  assign _01323_ = _01322_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5048" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[121];
  assign _01324_ = _01323_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5048" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[122];
  assign _01325_ = _01324_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5049" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[123];
  assign _01326_ = _01325_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5049" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[124];
  assign _01327_ = _01326_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5050" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[125];
  assign _01328_ = _01327_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5050" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[126];
  assign _01329_ = _01328_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5051" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[127];
  assign _01330_ = _01329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5051" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[128];
  assign _01331_ = _01330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5052" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[129];
  assign _01332_ = _01331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5052" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[130];
  assign _01333_ = _01332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5053" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[131];
  assign _01334_ = _01333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5053" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[132];
  assign _01335_ = _01334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5054" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[133];
  assign _01336_ = _01335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5054" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[134];
  assign _01337_ = _01336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5055" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[135];
  assign _01338_ = _01337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5055" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[136];
  assign _01339_ = _01338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5056" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[137];
  assign _01340_ = _01339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5056" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[138];
  assign _01341_ = _01340_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5057" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[139];
  assign _01342_ = _01341_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5057" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[140];
  assign _01343_ = _01342_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5058" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[141];
  assign _01344_ = _01343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5058" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[142];
  assign _01345_ = _01344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5059" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[143];
  assign _01346_ = _01345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5059" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[144];
  assign _01347_ = _01346_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5060" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[145];
  assign _01348_ = _01347_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5060" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[146];
  assign _01349_ = _01348_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5061" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[147];
  assign _01350_ = _01349_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5061" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[148];
  assign _01351_ = _01350_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5062" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[149];
  assign _01352_ = _01351_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5062" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[150];
  assign _01353_ = _01352_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5063" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[151];
  assign _01354_ = _01353_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5063" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[152];
  assign _01355_ = _01354_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5064" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[153];
  assign _01356_ = _01355_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5064" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[154];
  assign _01357_ = _01356_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5065" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[155];
  assign _01358_ = _01357_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5065" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[156];
  assign _01359_ = _01358_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5066" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[157];
  assign _01360_ = _01359_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5066" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[158];
  assign _01361_ = _01360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5067" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[159];
  assign _01362_ = _01361_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5067" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[160];
  assign _01363_ = _01362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5068" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[161];
  assign _01364_ = _01363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5068" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[162];
  assign _01365_ = _01364_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5069" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[163];
  assign _01366_ = _01365_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5069" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[164];
  assign _01367_ = _01366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5070" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[165];
  assign _01368_ = _01367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5070" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[166];
  assign _01369_ = _01368_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5071" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[167];
  assign _01370_ = _01369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5071" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[168];
  assign _01371_ = _01370_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5072" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[169];
  assign _01372_ = _01371_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5072" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[170];
  assign _01373_ = _01372_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5073" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[171];
  assign _01374_ = _01373_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5073" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[172];
  assign _01375_ = _01374_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5074" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[173];
  assign _01376_ = _01375_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5074" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[174];
  assign _01377_ = _01376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5075" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[175];
  assign _01378_ = _01377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5075" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[176];
  assign _01379_ = _01378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5076" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[177];
  assign _01380_ = _01379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5076" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[178];
  assign _01381_ = _01380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5077" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[179];
  assign _01382_ = _01381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5077" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[180];
  assign _01383_ = _01382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5078" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[181];
  assign _01384_ = _01383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5078" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[182];
  assign _01385_ = _01384_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5079" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[183];
  assign _01386_ = _01385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5079" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[184];
  assign _01387_ = _01386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5080" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[185];
  assign _01388_ = _01387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5080" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[186];
  assign _01389_ = _01388_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5081" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[187];
  assign _01390_ = _01389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5081" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[188];
  assign _01391_ = _01390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5082" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[189];
  assign _01392_ = _01391_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5082" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[190];
  assign _01393_ = _01392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5083" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[191];
  assign _01394_ = _01393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5083" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[192];
  assign _01395_ = _01394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5084" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[193];
  assign _01396_ = _01395_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5084" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[194];
  assign _01397_ = _01396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5085" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[195];
  assign _01398_ = _01397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5085" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[196];
  assign _01399_ = _01398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5086" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[197];
  assign _01400_ = _01399_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5086" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[198];
  assign _01401_ = _01400_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5087" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[199];
  assign _01402_ = _01401_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5087" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[200];
  assign _01403_ = _01402_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5088" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[201];
  assign _01404_ = _01403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5088" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[202];
  assign _01405_ = _01404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5089" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[203];
  assign _01406_ = _01405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5089" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[204];
  assign _01407_ = _01406_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5090" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[205];
  assign _01408_ = _01407_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5090" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[206];
  assign _01409_ = _01408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5091" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[207];
  assign _01410_ = _01409_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5091" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[208];
  assign _01411_ = _01410_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5092" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[209];
  assign _01412_ = _01411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5092" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[210];
  assign _01413_ = _01412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5093" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[211];
  assign _01414_ = _01413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5093" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[212];
  assign _01415_ = _01414_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5094" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[213];
  assign _01416_ = _01415_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5094" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[214];
  assign _01417_ = _01416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5095" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[215];
  assign _01418_ = _01417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5095" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[216];
  assign _01419_ = _01418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5096" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[217];
  assign _01420_ = _01419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5096" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[218];
  assign _01421_ = _01420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5097" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[219];
  assign _01422_ = _01421_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5097" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[220];
  assign _01423_ = _01422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5098" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[221];
  assign _01424_ = _01423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5098" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[222];
  assign _01425_ = _01424_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5099" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[223];
  assign _01426_ = _01425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5099" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[224];
  assign _01427_ = _01426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5100" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[225];
  assign _01428_ = _01427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5100" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[226];
  assign _01429_ = _01428_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5101" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[227];
  assign _01430_ = _01429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5101" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[228];
  assign _01431_ = _01430_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5102" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[229];
  assign _01432_ = _01431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5102" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[230];
  assign _01433_ = _01432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5103" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[231];
  assign _01434_ = _01433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5103" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[232];
  assign _01435_ = _01434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5104" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[233];
  assign _01436_ = _01435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5104" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[234];
  assign _01437_ = _01436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5105" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[235];
  assign _01438_ = _01437_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5105" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[236];
  assign _01439_ = _01438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5106" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[237];
  assign _01440_ = _01439_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5106" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[238];
  assign _01441_ = _01440_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5107" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[239];
  assign _01442_ = _01441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5107" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[240];
  assign _01443_ = _01442_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5108" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[241];
  assign _01444_ = _01443_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5108" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[242];
  assign _01445_ = _01444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5109" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[243];
  assign _01446_ = _01445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5109" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[244];
  assign _01447_ = _01446_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5110" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[245];
  assign _01448_ = _01447_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5110" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[246];
  assign _01449_ = _01448_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5111" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[247];
  assign _01450_ = _01449_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5111" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[248];
  assign _01451_ = _01450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5112" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[249];
  assign _01452_ = _01451_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5112" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[250];
  assign _01453_ = _01452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5113" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[251];
  assign _01454_ = _01453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5113" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[252];
  assign _01455_ = _01454_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5114" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[253];
  assign _01456_ = _01455_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5114" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[254];
  assign _01457_ = _01456_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5115" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[255];
  assign _01458_ = _01457_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5115" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[256];
  assign _01459_ = _01458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5116" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[257];
  assign _01460_ = _01459_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5116" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[258];
  assign _01461_ = _01460_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5117" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[259];
  assign _01462_ = _01461_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5117" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[260];
  assign _01463_ = _01462_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5118" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[261];
  assign _01464_ = _01463_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5118" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[262];
  assign _01465_ = _01464_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5119" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[263];
  assign _01466_ = _01465_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5119" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[264];
  assign _01467_ = _01466_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5120" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[265];
  assign _01468_ = _01467_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5120" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[266];
  assign _01469_ = _01468_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5121" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[267];
  assign _01470_ = _01469_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5121" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[268];
  assign _01471_ = _01470_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5122" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[269];
  assign _01472_ = _01471_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5122" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[270];
  assign _01473_ = _01472_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5123" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[271];
  assign _01474_ = _01473_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5123" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[272];
  assign _01475_ = _01474_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5124" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[273];
  assign _01476_ = _01475_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5124" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[274];
  assign _01477_ = _01476_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5125" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[275];
  assign _01478_ = _01477_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5125" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[276];
  assign _01479_ = _01478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5126" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[277];
  assign _01480_ = _01479_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5126" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[278];
  assign _01481_ = _01480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5127" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[279];
  assign _01482_ = _01481_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5127" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[280];
  assign _01483_ = _01482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5128" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[281];
  assign _01484_ = _01483_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5128" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[282];
  assign _01485_ = _01484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5129" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[283];
  assign _01486_ = _01485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5129" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[284];
  assign _01487_ = _01486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5130" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[285];
  assign _01488_ = _01487_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5130" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[286];
  assign _01489_ = _01488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5131" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[287];
  assign _01490_ = _01489_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5131" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[288];
  assign _01491_ = _01490_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5132" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[289];
  assign _01492_ = _01491_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5132" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[290];
  assign _01493_ = _01492_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5133" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[291];
  assign _01494_ = _01493_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5133" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[292];
  assign _01495_ = _01494_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5134" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[293];
  assign _01496_ = _01495_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5134" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[294];
  assign _01497_ = _01496_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5135" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[295];
  assign _01498_ = _01497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5135" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[296];
  assign _01499_ = _01498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5136" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[297];
  assign _01500_ = _01499_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5136" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[298];
  assign _01501_ = _01500_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5137" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[299];
  assign _01502_ = _01501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5137" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[300];
  assign _01503_ = _01502_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5138" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[301];
  assign _01504_ = _01503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5138" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[302];
  assign _01505_ = _01504_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5139" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[303];
  assign _01506_ = _01505_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5139" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[304];
  assign _01507_ = _01506_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5140" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[305];
  assign _01508_ = _01507_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5140" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[306];
  assign _01509_ = _01508_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5141" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[307];
  assign _01510_ = _01509_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5141" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[308];
  assign _01511_ = _01510_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5142" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[309];
  assign _01512_ = _01511_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5142" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[310];
  assign _01513_ = _01512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5143" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[311];
  assign _01514_ = _01513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5143" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[312];
  assign _01515_ = _01514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5144" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[313];
  assign _01516_ = _01515_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5144" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[314];
  assign _01517_ = _01516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5145" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[315];
  assign _01518_ = _01517_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5145" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[316];
  assign _01519_ = _01518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5146" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[317];
  assign _01520_ = _01519_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5146" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[318];
  assign _01521_ = _01520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5147" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[319];
  assign _01522_ = _01521_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5147" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[320];
  assign _01523_ = _01522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5148" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[321];
  assign _01524_ = _01523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5148" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[322];
  assign _01525_ = _01524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5149" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[323];
  assign _01526_ = _01525_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5149" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[324];
  assign _01527_ = _01526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5150" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[325];
  assign _01528_ = _01527_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5150" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[326];
  assign _01529_ = _01528_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5151" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[327];
  assign _01530_ = _01529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5151" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[328];
  assign _01531_ = _01530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5152" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[329];
  assign _01532_ = _01531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5152" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[330];
  assign _01533_ = _01532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5153" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[331];
  assign _01534_ = _01533_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5153" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[332];
  assign _01535_ = _01534_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5154" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[333];
  assign _01536_ = _01535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5154" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[334];
  assign _01537_ = _01536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5155" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[335];
  assign _01538_ = _01537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5155" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[336];
  assign _01539_ = _01538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5156" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[337];
  assign _01540_ = _01539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5156" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[338];
  assign _01541_ = _01540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5157" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[339];
  assign _01542_ = _01541_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5157" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[340];
  assign _01543_ = _01542_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5158" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[341];
  assign _01544_ = _01543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5158" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[342];
  assign _01545_ = _01544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5159" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[343];
  assign _01546_ = _01545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5159" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[344];
  assign _01547_ = _01546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5160" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[345];
  assign _01548_ = _01547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5160" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[346];
  assign _01549_ = _01548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5161" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[347];
  assign _01550_ = _01549_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5161" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[348];
  assign _01551_ = _01550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5162" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[349];
  assign _01552_ = _01551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5162" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[350];
  assign _01553_ = _01552_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5163" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[351];
  assign _01554_ = _01553_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5163" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[352];
  assign _01555_ = _01554_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5164" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[353];
  assign _01556_ = _01555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5164" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[354];
  assign _01557_ = _01556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5165" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[355];
  assign _01558_ = _01557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5165" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[356];
  assign _01559_ = _01558_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5166" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[357];
  assign _01560_ = _01559_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5166" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[358];
  assign _01561_ = _01560_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5167" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[359];
  assign _01562_ = _01561_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5167" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[360];
  assign _01563_ = _01562_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5168" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[361];
  assign _01564_ = _01563_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5168" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[362];
  assign _01565_ = _01564_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5169" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[363];
  assign _01566_ = _01565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5169" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[364];
  assign _01567_ = _01566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5170" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[365];
  assign _01568_ = _01567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5170" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[366];
  assign _01569_ = _01568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5171" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[367];
  assign _01570_ = _01569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5171" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[368];
  assign _01571_ = _01570_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5172" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[369];
  assign _01572_ = _01571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5172" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[370];
  assign _01573_ = _01572_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5173" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[371];
  assign _01574_ = _01573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5173" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[372];
  assign _01575_ = _01574_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5174" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[373];
  assign _01576_ = _01575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5174" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[374];
  assign _01577_ = _01576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5175" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[375];
  assign _01578_ = _01577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5175" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[376];
  assign _01579_ = _01578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5176" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[377];
  assign _01580_ = _01579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5176" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[378];
  assign _01581_ = _01580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5177" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[379];
  assign _01582_ = _01581_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5177" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[380];
  assign _01583_ = _01582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5178" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[381];
  assign _01584_ = _01583_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5178" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[382];
  assign _01585_ = _01584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5179" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[383];
  assign _01586_ = _01585_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5179" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[384];
  assign _01587_ = _01586_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5180" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[385];
  assign _01588_ = _01587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5180" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[386];
  assign _01589_ = _01588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5181" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[387];
  assign _01590_ = _01589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5181" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[388];
  assign _01591_ = _01590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5182" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[389];
  assign _01592_ = _01591_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5182" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[390];
  assign _01593_ = _01592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5183" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[391];
  assign _01594_ = _01593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5183" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[392];
  assign _01595_ = _01594_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5184" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[393];
  assign _01596_ = _01595_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5184" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[394];
  assign _01597_ = _01596_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5185" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[395];
  assign _01598_ = _01597_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5185" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[396];
  assign _01599_ = _01598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5186" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[397];
  assign _01600_ = _01599_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5186" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[398];
  assign _01601_ = _01600_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5187" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[399];
  assign _01602_ = _01601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5187" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[400];
  assign _01603_ = _01602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5188" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[401];
  assign _01604_ = _01603_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5188" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[402];
  assign _01605_ = _01604_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5189" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[403];
  assign _01606_ = _01605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5189" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[404];
  assign _01607_ = _01606_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5190" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[405];
  assign _01608_ = _01607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5190" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[406];
  assign _01609_ = _01608_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5191" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[407];
  assign _01610_ = _01609_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5191" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[408];
  assign _01611_ = _01610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5192" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[409];
  assign _01612_ = _01611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5192" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[410];
  assign _01613_ = _01612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5193" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[411];
  assign _01614_ = _01613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5193" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[412];
  assign _01615_ = _01614_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5194" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[413];
  assign _01616_ = _01615_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5194" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[414];
  assign _01617_ = _01616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5195" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[415];
  assign _01618_ = _01617_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5195" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[416];
  assign _01619_ = _01618_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5196" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[417];
  assign _01620_ = _01619_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5196" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[418];
  assign _01621_ = _01620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5197" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[419];
  assign _01622_ = _01621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5197" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[420];
  assign _01623_ = _01622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5198" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[421];
  assign _01624_ = _01623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5198" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[422];
  assign _01625_ = _01624_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5199" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[423];
  assign _01626_ = _01625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5199" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[424];
  assign _01627_ = _01626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5200" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[425];
  assign _01628_ = _01627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5200" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[426];
  assign _01629_ = _01628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5201" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[427];
  assign _01630_ = _01629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5201" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[428];
  assign _01631_ = _01630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5202" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[429];
  assign _01632_ = _01631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5202" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[430];
  assign _01633_ = _01632_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5203" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[431];
  assign _01634_ = _01633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5203" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[432];
  assign _01635_ = _01634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5204" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[433];
  assign _01636_ = _01635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5204" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[434];
  assign _01637_ = _01636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5205" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[435];
  assign _01638_ = _01637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5205" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[436];
  assign _01639_ = _01638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5206" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[437];
  assign _01640_ = _01639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5206" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[438];
  assign _01641_ = _01640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5207" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[439];
  assign _01642_ = _01641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5207" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[440];
  assign _01643_ = _01642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5208" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[441];
  assign _01644_ = _01643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5208" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[442];
  assign _01645_ = _01644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5209" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[443];
  assign _01646_ = _01645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5209" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[444];
  assign _01647_ = _01646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5210" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[445];
  assign _01648_ = _01647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5210" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[446];
  assign _01649_ = _01648_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5211" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[447];
  assign _01650_ = _01649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5211" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[448];
  assign _01651_ = _01650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5212" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[449];
  assign _01652_ = _01651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5212" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[450];
  assign _01653_ = _01652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5213" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[451];
  assign _01654_ = _01653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5213" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[452];
  assign _01655_ = _01654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5214" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[453];
  assign _01656_ = _01655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5214" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[454];
  assign _01657_ = _01656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5215" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[455];
  assign _01658_ = _01657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5215" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[456];
  assign _01659_ = _01658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5216" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[457];
  assign _01660_ = _01659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5216" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[458];
  assign _01661_ = _01660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5217" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[459];
  assign _01662_ = _01661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5217" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[460];
  assign _01663_ = _01662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5218" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[461];
  assign _01664_ = _01663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5218" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[462];
  assign _01665_ = _01664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5219" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[463];
  assign _01666_ = _01665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5219" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[464];
  assign _01667_ = _01666_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5220" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[465];
  assign _01668_ = _01667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5220" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[466];
  assign _01669_ = _01668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5221" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[467];
  assign _01670_ = _01669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5221" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[468];
  assign _01671_ = _01670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5222" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[469];
  assign _01672_ = _01671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5222" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[470];
  assign _01673_ = _01672_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5223" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[471];
  assign _01674_ = _01673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5223" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[472];
  assign _01675_ = _01674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5224" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[473];
  assign _01676_ = _01675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5224" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[474];
  assign _01677_ = _01676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5225" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[475];
  assign _01678_ = _01677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5225" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[476];
  assign _01679_ = _01678_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5226" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[477];
  assign _01680_ = _01679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5226" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[478];
  assign _01681_ = _01680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5227" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[479];
  assign _01682_ = _01681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5227" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[480];
  assign _01683_ = _01682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5228" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[481];
  assign _01684_ = _01683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5228" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[482];
  assign _01685_ = _01684_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5229" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[483];
  assign _01686_ = _01685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5229" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[484];
  assign _01687_ = _01686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5230" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[485];
  assign _01688_ = _01687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5230" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[486];
  assign _01689_ = _01688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5231" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[487];
  assign _01690_ = _01689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5231" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[488];
  assign _01691_ = _01690_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5232" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[489];
  assign _01692_ = _01691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5232" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[490];
  assign _01693_ = _01692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5233" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[491];
  assign _01694_ = _01693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5233" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[492];
  assign _01695_ = _01694_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5234" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[493];
  assign _01696_ = _01695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5234" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[494];
  assign _01697_ = _01696_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5235" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[495];
  assign _01698_ = _01697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5235" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[496];
  assign _01699_ = _01698_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5236" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[497];
  assign _01700_ = _01699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5236" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[498];
  assign _01701_ = _01700_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5237" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[499];
  assign _01702_ = _01701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5237" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[500];
  assign _01703_ = _01702_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5238" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[501];
  assign _01704_ = _01703_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5238" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[502];
  assign _01705_ = _01704_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5239" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[503];
  assign _01706_ = _01705_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5239" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[504];
  assign _01707_ = _01706_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5240" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[505];
  assign _01708_ = _01707_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5240" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[506];
  assign _01709_ = _01708_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5241" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[507];
  assign _01710_ = _01709_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5241" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[508];
  assign _01711_ = _01710_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5242" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[509];
  assign _01712_ = _01711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5242" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[510];
  assign _01713_ = _01712_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5243" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[511];
  assign _01714_ = _01713_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5243" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[512];
  assign _01715_ = _01714_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5244" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[513];
  assign _01716_ = _01715_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5244" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[514];
  assign _01717_ = _01716_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5245" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[515];
  assign _01718_ = _01717_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5245" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[516];
  assign _01719_ = _01718_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5246" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[517];
  assign _01720_ = _01719_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5246" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[518];
  assign _01721_ = _01720_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5247" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[519];
  assign _01722_ = _01721_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5247" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[520];
  assign _01723_ = _01722_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5248" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[521];
  assign _01724_ = _01723_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5248" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[522];
  assign _01725_ = _01724_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5249" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[523];
  assign _01726_ = _01725_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5249" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[524];
  assign _01727_ = _01726_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5250" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[525];
  assign _01728_ = _01727_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5250" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[526];
  assign _01729_ = _01728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5251" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[527];
  assign _01730_ = _01729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5251" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[528];
  assign _01731_ = _01730_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5252" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[529];
  assign _01732_ = _01731_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5252" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[530];
  assign _01733_ = _01732_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5253" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[531];
  assign _01734_ = _01733_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5253" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[532];
  assign _01735_ = _01734_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5254" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[533];
  assign _01736_ = _01735_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5254" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[534];
  assign _01737_ = _01736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5255" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[535];
  assign _01738_ = _01737_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5255" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[536];
  assign _01739_ = _01738_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5256" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[537];
  assign _01740_ = _01739_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5256" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[538];
  assign _01741_ = _01740_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5257" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[539];
  assign _01742_ = _01741_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5257" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[540];
  assign _01743_ = _01742_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5258" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[541];
  assign _01744_ = _01743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5258" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[542];
  assign _01745_ = _01744_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5259" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[543];
  assign _01746_ = _01745_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5259" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[544];
  assign _01747_ = _01746_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5260" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[545];
  assign _01748_ = _01747_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5260" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[546];
  assign _01749_ = _01748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5261" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[547];
  assign _01750_ = _01749_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5261" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[548];
  assign _01751_ = _01750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5262" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[549];
  assign _01752_ = _01751_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5262" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[550];
  assign _01753_ = _01752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5263" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[551];
  assign _01754_ = _01753_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5263" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[552];
  assign _01755_ = _01754_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5264" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[553];
  assign _01756_ = _01755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5264" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[554];
  assign _01757_ = _01756_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5265" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[555];
  assign _01758_ = _01757_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5265" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[556];
  assign _01759_ = _01758_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5266" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[557];
  assign _01760_ = _01759_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5266" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[558];
  assign _01761_ = _01760_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5267" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[559];
  assign _01762_ = _01761_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5267" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[560];
  assign _01763_ = _01762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5268" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[561];
  assign _01764_ = _01763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5268" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[562];
  assign _01765_ = _01764_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5269" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[563];
  assign _01766_ = _01765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5269" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[564];
  assign _01767_ = _01766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5270" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[565];
  assign _01768_ = _01767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5270" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[566];
  assign _01769_ = _01768_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5271" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[567];
  assign _01770_ = _01769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5271" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[568];
  assign _01771_ = _01770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5272" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[569];
  assign _01772_ = _01771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5272" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[570];
  assign _01773_ = _01772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5273" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[571];
  assign _01774_ = _01773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5273" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[572];
  assign _01775_ = _01774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5274" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[573];
  assign _01776_ = _01775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5274" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[574];
  assign _01777_ = _01776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5275" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[575];
  assign _01778_ = _01777_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5275" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[576];
  assign _01779_ = _01778_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5276" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[577];
  assign _01780_ = _01779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5276" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[578];
  assign _01781_ = _01780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5277" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[579];
  assign _01782_ = _01781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5277" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[580];
  assign _01783_ = _01782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5278" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[581];
  assign _01784_ = _01783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5278" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[582];
  assign _01785_ = _01784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5279" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[583];
  assign _01786_ = _01785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5279" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[584];
  assign _01787_ = _01786_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5280" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[585];
  assign _01788_ = _01787_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5280" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[586];
  assign _01789_ = _01788_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5281" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[587];
  assign _01790_ = _01789_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5281" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[588];
  assign _01791_ = _01790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5282" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[589];
  assign _01792_ = _01791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5282" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[590];
  assign _01793_ = _01792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5283" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[591];
  assign _01794_ = _01793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5283" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[592];
  assign _01795_ = _01794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5284" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[593];
  assign _01796_ = _01795_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5284" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[594];
  assign _01797_ = _01796_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5285" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[595];
  assign _01798_ = _01797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5285" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[596];
  assign _01799_ = _01798_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5286" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[597];
  assign _01800_ = _01799_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5286" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[598];
  assign _01801_ = _01800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5287" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[599];
  assign _01802_ = _01801_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5287" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[600];
  assign _01803_ = _01802_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5288" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[601];
  assign _01804_ = _01803_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5288" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[602];
  assign _01805_ = _01804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5289" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[603];
  assign _01806_ = _01805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5289" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[604];
  assign _01807_ = _01806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5290" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[605];
  assign _01808_ = _01807_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5290" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[606];
  assign _01809_ = _01808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5291" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[607];
  assign _01810_ = _01809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5291" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[608];
  assign _01811_ = _01810_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5292" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[609];
  assign _01812_ = _01811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5292" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[610];
  assign _01813_ = _01812_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5293" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[611];
  assign _01814_ = _01813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5293" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[612];
  assign _01815_ = _01814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5294" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[613];
  assign _01816_ = _01815_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5294" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[614];
  assign _01817_ = _01816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5295" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[615];
  assign _01818_ = _01817_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5295" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[616];
  assign _01819_ = _01818_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5296" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[617];
  assign _01820_ = _01819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5296" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[618];
  assign _01821_ = _01820_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5297" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[619];
  assign _01822_ = _01821_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5297" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[620];
  assign _01823_ = _01822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5298" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[621];
  assign _01824_ = _01823_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5298" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[622];
  assign _01825_ = _01824_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5299" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[623];
  assign _01826_ = _01825_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5299" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[624];
  assign _01827_ = _01826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5300" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[625];
  assign _01828_ = _01827_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5300" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[626];
  assign _01829_ = _01828_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5301" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[627];
  assign _01830_ = _01829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5301" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[628];
  assign _01831_ = _01830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5302" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[629];
  assign _01832_ = _01831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5302" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[630];
  assign _01833_ = _01832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5303" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[631];
  assign _01834_ = _01833_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5303" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[632];
  assign _01835_ = _01834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5304" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[633];
  assign _01836_ = _01835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5304" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[634];
  assign _01837_ = _01836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5305" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[635];
  assign _01838_ = _01837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5305" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[636];
  assign _01839_ = _01838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5306" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[637];
  assign _01840_ = _01839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5306" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[638];
  assign _01841_ = _01840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5307" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[639];
  assign _01842_ = _01841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5307" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[640];
  assign _01843_ = _01842_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5308" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[641];
  assign _01844_ = _01843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5308" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[642];
  assign _01845_ = _01844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5309" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[643];
  assign _01846_ = _01845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5309" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[644];
  assign _01847_ = _01846_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5310" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[645];
  assign _01848_ = _01847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5310" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[646];
  assign _01849_ = _01848_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5311" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[647];
  assign _01850_ = _01849_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5311" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[648];
  assign _01851_ = _01850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5312" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[649];
  assign _01852_ = _01851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5312" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[650];
  assign _01853_ = _01852_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5313" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[651];
  assign _01854_ = _01853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5313" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[652];
  assign _01855_ = _01854_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5314" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[653];
  assign _01856_ = _01855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5314" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[654];
  assign _01857_ = _01856_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5315" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[655];
  assign _01858_ = _01857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5315" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[656];
  assign _01859_ = _01858_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5316" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[657];
  assign _01860_ = _01859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5316" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[658];
  assign _01861_ = _01860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5317" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[659];
  assign _01862_ = _01861_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5317" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[660];
  assign _01863_ = _01862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5318" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[661];
  assign _01864_ = _01863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5318" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[662];
  assign _01865_ = _01864_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5319" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[663];
  assign _01866_ = _01865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5319" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[664];
  assign _01867_ = _01866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5320" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[665];
  assign _01868_ = _01867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5320" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[666];
  assign _01869_ = _01868_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5321" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[667];
  assign _01870_ = _01869_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5321" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[668];
  assign _01871_ = _01870_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5322" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[669];
  assign _01872_ = _01871_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5322" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[670];
  assign _01873_ = _01872_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5323" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[671];
  assign _01874_ = _01873_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5323" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[672];
  assign _01875_ = _01874_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5324" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[673];
  assign _01876_ = _01875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5324" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[674];
  assign _01877_ = _01876_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5325" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[675];
  assign _01878_ = _01877_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5325" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[676];
  assign _01879_ = _01878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5326" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[677];
  assign _01880_ = _01879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5326" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[678];
  assign _01881_ = _01880_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5327" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[679];
  assign _01882_ = _01881_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5327" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[680];
  assign _01883_ = _01882_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5328" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[681];
  assign _01884_ = _01883_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5328" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[682];
  assign _01885_ = _01884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5329" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[683];
  assign _01886_ = _01885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5329" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[684];
  assign _01887_ = _01886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5330" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[685];
  assign _01888_ = _01887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5330" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[686];
  assign _01889_ = _01888_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5331" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[687];
  assign _01890_ = _01889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5331" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[688];
  assign _01891_ = _01890_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5332" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[689];
  assign _01892_ = _01891_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5332" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[690];
  assign _01893_ = _01892_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5333" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[691];
  assign _01894_ = _01893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5333" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[692];
  assign _01895_ = _01894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5334" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[693];
  assign _01896_ = _01895_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5334" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[694];
  assign _01897_ = _01896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5335" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[695];
  assign _01898_ = _01897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5335" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[696];
  assign _01899_ = _01898_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5336" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[697];
  assign _01900_ = _01899_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5336" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[698];
  assign _01901_ = _01900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5337" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[699];
  assign _01902_ = _01901_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5337" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[700];
  assign _01903_ = _01902_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5338" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[701];
  assign _01904_ = _01903_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5338" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[702];
  assign _01905_ = _01904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5339" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[703];
  assign _01906_ = _01905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5339" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[704];
  assign _01907_ = _01906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5340" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[705];
  assign _01908_ = _01907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5340" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[706];
  assign _01909_ = _01908_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5341" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[707];
  assign _01910_ = _01909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5341" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[708];
  assign _01911_ = _01910_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5342" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[709];
  assign _01912_ = _01911_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5342" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[710];
  assign _01913_ = _01912_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5343" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[711];
  assign _01914_ = _01913_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5343" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[712];
  assign _01915_ = _01914_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5344" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[713];
  assign _01916_ = _01915_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5344" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[714];
  assign _01917_ = _01916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5345" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[715];
  assign _01918_ = _01917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5345" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[716];
  assign _01919_ = _01918_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5346" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[717];
  assign _01920_ = _01919_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5346" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[718];
  assign _01921_ = _01920_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5347" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[719];
  assign _01922_ = _01921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5347" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[720];
  assign _01923_ = _01922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5348" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[721];
  assign _01924_ = _01923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5348" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[722];
  assign _01925_ = _01924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5349" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[723];
  assign _01926_ = _01925_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5349" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[724];
  assign _01927_ = _01926_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5350" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[725];
  assign _01928_ = _01927_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5350" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[726];
  assign _01929_ = _01928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5351" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[727];
  assign _01930_ = _01929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5351" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[728];
  assign _01931_ = _01930_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5352" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[729];
  assign _01932_ = _01931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5352" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[730];
  assign _01933_ = _01932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5353" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[731];
  assign _01934_ = _01933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5353" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[732];
  assign _01935_ = _01934_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5354" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[733];
  assign _01936_ = _01935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5354" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[734];
  assign _01937_ = _01936_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5355" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[735];
  assign _01938_ = _01937_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5355" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[736];
  assign _01939_ = _01938_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5356" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[737];
  assign _01940_ = _01939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5356" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[738];
  assign _01941_ = _01940_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5357" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[739];
  assign _01942_ = _01941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5357" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[740];
  assign _01943_ = _01942_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5358" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[741];
  assign _01944_ = _01943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5358" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[742];
  assign _01945_ = _01944_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5359" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[743];
  assign _01946_ = _01945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5359" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[744];
  assign _01947_ = _01946_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5360" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[745];
  assign _01948_ = _01947_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5360" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[746];
  assign _01949_ = _01948_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5361" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[747];
  assign _01950_ = _01949_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5361" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[748];
  assign _01951_ = _01950_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5362" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[749];
  assign _01952_ = _01951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5362" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[750];
  assign _01953_ = _01952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5363" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[751];
  assign _01954_ = _01953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5363" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[752];
  assign _01955_ = _01954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5364" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[753];
  assign _01956_ = _01955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5364" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[754];
  assign _01957_ = _01956_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5365" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[755];
  assign _01958_ = _01957_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5365" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[756];
  assign _01959_ = _01958_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5366" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[757];
  assign _01960_ = _01959_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5366" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[758];
  assign _01961_ = _01960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5367" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[759];
  assign _01962_ = _01961_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5367" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[760];
  assign _01963_ = _01962_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5368" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[761];
  assign _01964_ = _01963_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5368" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[762];
  assign _01965_ = _01964_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5369" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[763];
  assign _01966_ = _01965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5369" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[764];
  assign _01967_ = _01966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5370" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[765];
  assign _01968_ = _01967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5370" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[766];
  assign _01969_ = _01968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5371" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[767];
  assign _01970_ = _01969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5371" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[768];
  assign _01971_ = _01970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5372" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[769];
  assign _01972_ = _01971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5372" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[770];
  assign _01973_ = _01972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5373" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[771];
  assign _01974_ = _01973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5373" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[772];
  assign _01975_ = _01974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5374" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[773];
  assign _01976_ = _01975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5374" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[774];
  assign _01977_ = _01976_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5375" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[775];
  assign _01978_ = _01977_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5375" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[776];
  assign _01979_ = _01978_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5376" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[777];
  assign _01980_ = _01979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5376" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[778];
  assign _01981_ = _01980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5377" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[779];
  assign _01982_ = _01981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5377" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[780];
  assign _01983_ = _01982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5378" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[781];
  assign _01984_ = _01983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5378" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[782];
  assign _01985_ = _01984_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5379" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[783];
  assign _01986_ = _01985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5379" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[784];
  assign _01987_ = _01986_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5380" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[785];
  assign _01988_ = _01987_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5380" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[786];
  assign _01989_ = _01988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5381" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[787];
  assign _01990_ = _01989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5381" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[788];
  assign _01991_ = _01990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5382" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[789];
  assign _01992_ = _01991_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5382" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[790];
  assign _01993_ = _01992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5383" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[791];
  assign _01994_ = _01993_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5383" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[792];
  assign _01995_ = _01994_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5384" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[793];
  assign _01996_ = _01995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5384" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[794];
  assign _01997_ = _01996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5385" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[795];
  assign _01998_ = _01997_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5385" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[796];
  assign _01999_ = _01998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5386" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[797];
  assign _02000_ = _01999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5386" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[798];
  assign _02001_ = _02000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5387" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[799];
  assign _02002_ = _02001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5387" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[800];
  assign _02003_ = _02002_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5388" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[801];
  assign _02004_ = _02003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5388" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[802];
  assign _02005_ = _02004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5389" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[803];
  assign _02006_ = _02005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5389" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[804];
  assign _02007_ = _02006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5390" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[805];
  assign _02008_ = _02007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5390" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[806];
  assign _02009_ = _02008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5391" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[807];
  assign _02010_ = _02009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5391" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[808];
  assign _02011_ = _02010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5392" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[809];
  assign _02012_ = _02011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5392" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[810];
  assign _02013_ = _02012_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5393" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[811];
  assign _02014_ = _02013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5393" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[812];
  assign _02015_ = _02014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5394" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[813];
  assign _02016_ = _02015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5394" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[814];
  assign _02017_ = _02016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5395" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[815];
  assign _02018_ = _02017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5395" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[816];
  assign _02019_ = _02018_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5396" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[817];
  assign _02020_ = _02019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5396" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[818];
  assign _02021_ = _02020_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5397" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[819];
  assign _02022_ = _02021_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5397" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[820];
  assign _02023_ = _02022_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5398" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[821];
  assign _02024_ = _02023_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5398" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[822];
  assign _02025_ = _02024_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5399" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[823];
  assign _02026_ = _02025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5399" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[824];
  assign _02027_ = _02026_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5400" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[825];
  assign _02028_ = _02027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5400" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[826];
  assign _02029_ = _02028_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5401" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[827];
  assign _02030_ = _02029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5401" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[828];
  assign _02031_ = _02030_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5402" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[829];
  assign _02032_ = _02031_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5402" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[830];
  assign _02033_ = _02032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5403" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[831];
  assign _02034_ = _02033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5403" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[832];
  assign _02035_ = _02034_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5404" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[833];
  assign _02036_ = _02035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5404" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[834];
  assign _02037_ = _02036_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5405" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[835];
  assign _02038_ = _02037_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5405" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[836];
  assign _02039_ = _02038_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5406" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[837];
  assign _02040_ = _02039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5406" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[838];
  assign _02041_ = _02040_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5407" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[839];
  assign _02042_ = _02041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5407" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[840];
  assign _02043_ = _02042_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5408" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[841];
  assign _02044_ = _02043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5408" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[842];
  assign _02045_ = _02044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5409" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[843];
  assign _02046_ = _02045_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5409" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[844];
  assign _02047_ = _02046_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5410" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[845];
  assign _02048_ = _02047_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5410" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[846];
  assign _02049_ = _02048_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5411" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[847];
  assign _02050_ = _02049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5411" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[848];
  assign _02051_ = _02050_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5412" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[849];
  assign _02052_ = _02051_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5412" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[850];
  assign _02053_ = _02052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5413" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[851];
  assign _02054_ = _02053_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5413" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[852];
  assign _02055_ = _02054_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5414" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[853];
  assign _02056_ = _02055_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5414" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[854];
  assign _02057_ = _02056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5415" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[855];
  assign _02058_ = _02057_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5415" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[856];
  assign _02059_ = _02058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5416" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[857];
  assign _02060_ = _02059_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5416" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[858];
  assign _02061_ = _02060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5417" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[859];
  assign _02062_ = _02061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5417" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[860];
  assign _02063_ = _02062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5418" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[861];
  assign _02064_ = _02063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5418" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[862];
  assign _02065_ = _02064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5419" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[863];
  assign _02066_ = _02065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5419" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[864];
  assign _02067_ = _02066_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5420" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[865];
  assign _02068_ = _02067_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5420" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[866];
  assign _02069_ = _02068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5421" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[867];
  assign _02070_ = _02069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5421" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[868];
  assign _02071_ = _02070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5422" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[869];
  assign _02072_ = _02071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5422" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[870];
  assign _02073_ = _02072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5423" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[871];
  assign _02074_ = _02073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5423" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[872];
  assign _02075_ = _02074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5424" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[873];
  assign _02076_ = _02075_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5424" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[874];
  assign _02077_ = _02076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5425" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[875];
  assign _02078_ = _02077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5425" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[876];
  assign _02079_ = _02078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5426" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[877];
  assign _02080_ = _02079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5426" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[878];
  assign _02081_ = _02080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5427" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[879];
  assign _02082_ = _02081_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5427" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[880];
  assign _02083_ = _02082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5428" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[881];
  assign _02084_ = _02083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5428" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[882];
  assign _02085_ = _02084_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5429" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[883];
  assign _02086_ = _02085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5429" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[884];
  assign _02087_ = _02086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5430" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[885];
  assign _02088_ = _02087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5430" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[886];
  assign _02089_ = _02088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5431" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[887];
  assign _02090_ = _02089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5431" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[888];
  assign _02091_ = _02090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5432" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[889];
  assign _02092_ = _02091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5432" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[890];
  assign _02093_ = _02092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5433" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[891];
  assign _02094_ = _02093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5433" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[892];
  assign _02095_ = _02094_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5434" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[893];
  assign _02096_ = _02095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5434" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[894];
  assign _02097_ = _02096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5435" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[895];
  assign _02098_ = _02097_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5435" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[896];
  assign _02099_ = _02098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5436" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[897];
  assign _02100_ = _02099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5436" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[898];
  assign _02101_ = _02100_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5437" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[899];
  assign _02102_ = _02101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5437" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[900];
  assign _02103_ = _02102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5438" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[901];
  assign _02104_ = _02103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5438" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[902];
  assign _02105_ = _02104_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5439" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[903];
  assign _02106_ = _02105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5439" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[904];
  assign _02107_ = _02106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5440" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[905];
  assign _02108_ = _02107_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5440" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[906];
  assign _02109_ = _02108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5441" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[907];
  assign _02110_ = _02109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5441" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[908];
  assign _02111_ = _02110_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5442" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[909];
  assign _02112_ = _02111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5442" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[910];
  assign _02113_ = _02112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5443" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[911];
  assign _02114_ = _02113_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5443" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[912];
  assign _02115_ = _02114_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5444" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[913];
  assign _02116_ = _02115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5444" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[914];
  assign _02117_ = _02116_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5445" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[915];
  assign _02118_ = _02117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5445" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[916];
  assign _02119_ = _02118_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5446" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[917];
  assign _02120_ = _02119_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5446" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[918];
  assign _02121_ = _02120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5447" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[919];
  assign _02122_ = _02121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5447" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[920];
  assign _02123_ = _02122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5448" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[921];
  assign _02124_ = _02123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5448" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[922];
  assign _02125_ = _02124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5449" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[923];
  assign _02126_ = _02125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5449" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[924];
  assign _02127_ = _02126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5450" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[925];
  assign _02128_ = _02127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5450" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[926];
  assign _02129_ = _02128_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5451" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[927];
  assign _02130_ = _02129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5451" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[928];
  assign _02131_ = _02130_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5452" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[929];
  assign _02132_ = _02131_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5452" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[930];
  assign _02133_ = _02132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5453" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[931];
  assign _02134_ = _02133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5453" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[932];
  assign _02135_ = _02134_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5454" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[933];
  assign _02136_ = _02135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5454" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[934];
  assign _02137_ = _02136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5455" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[935];
  assign _02138_ = _02137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5455" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[936];
  assign _02139_ = _02138_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5456" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[937];
  assign _02140_ = _02139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5456" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[938];
  assign _02141_ = _02140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5457" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[939];
  assign _02142_ = _02141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5457" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[940];
  assign _02143_ = _02142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5458" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[941];
  assign _02144_ = _02143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5458" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[942];
  assign _02145_ = _02144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5459" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[943];
  assign _02146_ = _02145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5459" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[944];
  assign _02147_ = _02146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5460" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[945];
  assign _02148_ = _02147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5460" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[946];
  assign _02149_ = _02148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5461" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[947];
  assign _02150_ = _02149_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5461" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[948];
  assign _02151_ = _02150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5462" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[949];
  assign _02152_ = _02151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5462" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[950];
  assign _02153_ = _02152_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5463" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[951];
  assign _02154_ = _02153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5463" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[952];
  assign _02155_ = _02154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5464" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[953];
  assign _02156_ = _02155_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5464" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[954];
  assign _02157_ = _02156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5465" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[955];
  assign _02158_ = _02157_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5465" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[956];
  assign _02159_ = _02158_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5466" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[957];
  assign _02160_ = _02159_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5466" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[958];
  assign _02161_ = _02160_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5467" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[959];
  assign _02162_ = _02161_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5467" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[960];
  assign _02163_ = _02162_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5468" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[961];
  assign _02164_ = _02163_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5468" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[962];
  assign _02165_ = _02164_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5469" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[963];
  assign _02166_ = _02165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5469" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[964];
  assign _02167_ = _02166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5470" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[965];
  assign _02168_ = _02167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5470" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[966];
  assign _02169_ = _02168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5471" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[967];
  assign _02170_ = _02169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5471" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[968];
  assign _02171_ = _02170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5472" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[969];
  assign _02172_ = _02171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5472" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[970];
  assign _02173_ = _02172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5473" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[971];
  assign _02174_ = _02173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5473" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[972];
  assign _02175_ = _02174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5474" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[973];
  assign _02176_ = _02175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5474" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[974];
  assign _02177_ = _02176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5475" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[975];
  assign _02178_ = _02177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5475" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[976];
  assign _02179_ = _02178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5476" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[977];
  assign _02180_ = _02179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5476" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[978];
  assign _02181_ = _02180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5477" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[979];
  assign _02182_ = _02181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5477" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[980];
  assign _02183_ = _02182_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5478" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[981];
  assign _02184_ = _02183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5478" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[982];
  assign _02185_ = _02184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5479" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[983];
  assign _02186_ = _02185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5479" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[984];
  assign _02187_ = _02186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5480" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[985];
  assign _02188_ = _02187_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5480" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[986];
  assign _02189_ = _02188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5481" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[987];
  assign _02190_ = _02189_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5481" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[988];
  assign _02191_ = _02190_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5482" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[989];
  assign _02192_ = _02191_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5482" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[990];
  assign _02193_ = _02192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5483" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[991];
  assign _02194_ = _02193_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5483" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[992];
  assign _02195_ = _02194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5484" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[993];
  assign _02196_ = _02195_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5484" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[994];
  assign _02197_ = _02196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5485" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[995];
  assign _02198_ = _02197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5485" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[996];
  assign _02199_ = _02198_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5486" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[997];
  assign _02200_ = _02199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5486" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[998];
  assign _02201_ = _02200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5487" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[999];
  assign _02202_ = _02201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5487" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1000];
  assign _02203_ = _02202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5488" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1001];
  assign _02204_ = _02203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5488" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1002];
  assign _02205_ = _02204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5489" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1003];
  assign _02206_ = _02205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5489" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1004];
  assign _02207_ = _02206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5490" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1005];
  assign _02208_ = _02207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5490" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1006];
  assign _02209_ = _02208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5491" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1007];
  assign _02210_ = _02209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5491" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1008];
  assign _02211_ = _02210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5492" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1009];
  assign _02212_ = _02211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5492" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1010];
  assign _02213_ = _02212_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5493" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1011];
  assign _02214_ = _02213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5493" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1012];
  assign _02215_ = _02214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5494" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1013];
  assign _02216_ = _02215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5494" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1014];
  assign _02217_ = _02216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5495" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1015];
  assign _02218_ = _02217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5495" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1016];
  assign _02219_ = _02218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5496" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1017];
  assign _02220_ = _02219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5496" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1018];
  assign _02221_ = _02220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5497" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1019];
  assign _02222_ = _02221_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5497" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1020];
  assign _02223_ = _02222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5498" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva[1021];
  assign _02224_ = _02223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5498" *) _00854_;
  assign _02225_ = IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5504" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1];
  assign _02226_ = _02225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5504" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[2];
  assign _02227_ = _02226_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5505" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[3];
  assign _02228_ = _02227_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5505" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[4];
  assign _02229_ = _02228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5506" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[5];
  assign _02230_ = _02229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5506" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[6];
  assign _02231_ = _02230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5507" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[7];
  assign _02232_ = _02231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5507" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[8];
  assign _02233_ = _02232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5508" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[9];
  assign _02234_ = _02233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5508" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[10];
  assign _02235_ = _02234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5509" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[11];
  assign _02236_ = _02235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5509" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[12];
  assign _02237_ = _02236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5510" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[13];
  assign _02238_ = _02237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5510" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[14];
  assign _02239_ = _02238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5511" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[15];
  assign _02240_ = _02239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5511" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[16];
  assign _02241_ = _02240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5512" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[17];
  assign _02242_ = _02241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5512" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[18];
  assign _02243_ = _02242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5513" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[19];
  assign _02244_ = _02243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5513" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[20];
  assign _02245_ = _02244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5514" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[21];
  assign _02246_ = _02245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5514" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[22];
  assign _02247_ = _02246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5515" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[23];
  assign _02248_ = _02247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5515" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[24];
  assign _02249_ = _02248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5516" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[25];
  assign _02250_ = _02249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5516" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[26];
  assign _02251_ = _02250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5517" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[27];
  assign _02252_ = _02251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5517" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[28];
  assign _02253_ = _02252_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5518" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[29];
  assign _02254_ = _02253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5518" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[30];
  assign _02255_ = _02254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5519" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[31];
  assign _02256_ = _02255_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5519" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[32];
  assign _02257_ = _02256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5520" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[33];
  assign _02258_ = _02257_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5520" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[34];
  assign _02259_ = _02258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5521" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[35];
  assign _02260_ = _02259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5521" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[36];
  assign _02261_ = _02260_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5522" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[37];
  assign _02262_ = _02261_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5522" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[38];
  assign _02263_ = _02262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5523" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[39];
  assign _02264_ = _02263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5523" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[40];
  assign _02265_ = _02264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5524" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[41];
  assign _02266_ = _02265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5524" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[42];
  assign _02267_ = _02266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5525" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[43];
  assign _02268_ = _02267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5525" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[44];
  assign _02269_ = _02268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5526" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[45];
  assign _02270_ = _02269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5526" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[46];
  assign _02271_ = _02270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5527" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[47];
  assign _02272_ = _02271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5527" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[48];
  assign _02273_ = _02272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5528" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[49];
  assign _02274_ = _02273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5528" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[50];
  assign _02275_ = _02274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5529" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[51];
  assign _02276_ = _02275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5529" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[52];
  assign _02277_ = _02276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5530" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[53];
  assign _02278_ = _02277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5530" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[54];
  assign _02279_ = _02278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5531" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[55];
  assign _02280_ = _02279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5531" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[56];
  assign _02281_ = _02280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5532" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[57];
  assign _02282_ = _02281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5532" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[58];
  assign _02283_ = _02282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5533" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[59];
  assign _02284_ = _02283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5533" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[60];
  assign _02285_ = _02284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5534" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[61];
  assign _02286_ = _02285_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5534" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[62];
  assign _02287_ = _02286_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5535" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[63];
  assign _02288_ = _02287_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5535" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[64];
  assign _02289_ = _02288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5536" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[65];
  assign _02290_ = _02289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5536" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[66];
  assign _02291_ = _02290_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5537" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[67];
  assign _02292_ = _02291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5537" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[68];
  assign _02293_ = _02292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5538" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[69];
  assign _02294_ = _02293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5538" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[70];
  assign _02295_ = _02294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5539" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[71];
  assign _02296_ = _02295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5539" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[72];
  assign _02297_ = _02296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5540" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[73];
  assign _02298_ = _02297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5540" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[74];
  assign _02299_ = _02298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5541" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[75];
  assign _02300_ = _02299_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5541" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[76];
  assign _02301_ = _02300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5542" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[77];
  assign _02302_ = _02301_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5542" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[78];
  assign _02303_ = _02302_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5543" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[79];
  assign _02304_ = _02303_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5543" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[80];
  assign _02305_ = _02304_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5544" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[81];
  assign _02306_ = _02305_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5544" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[82];
  assign _02307_ = _02306_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5545" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[83];
  assign _02308_ = _02307_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5545" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[84];
  assign _02309_ = _02308_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5546" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[85];
  assign _02310_ = _02309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5546" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[86];
  assign _02311_ = _02310_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5547" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[87];
  assign _02312_ = _02311_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5547" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[88];
  assign _02313_ = _02312_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5548" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[89];
  assign _02314_ = _02313_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5548" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[90];
  assign _02315_ = _02314_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5549" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[91];
  assign _02316_ = _02315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5549" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[92];
  assign _02317_ = _02316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5550" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[93];
  assign _02318_ = _02317_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5550" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[94];
  assign _02319_ = _02318_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5551" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[95];
  assign _02320_ = _02319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5551" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[96];
  assign _02321_ = _02320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5552" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[97];
  assign _02322_ = _02321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5552" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[98];
  assign _02323_ = _02322_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5553" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[99];
  assign _02324_ = _02323_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5553" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[100];
  assign _02325_ = _02324_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5554" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[101];
  assign _02326_ = _02325_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5554" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[102];
  assign _02327_ = _02326_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5555" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[103];
  assign _02328_ = _02327_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5555" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[104];
  assign _02329_ = _02328_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5556" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[105];
  assign _02330_ = _02329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5556" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[106];
  assign _02331_ = _02330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5557" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[107];
  assign _02332_ = _02331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5557" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[108];
  assign _02333_ = _02332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5558" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[109];
  assign _02334_ = _02333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5558" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[110];
  assign _02335_ = _02334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5559" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[111];
  assign _02336_ = _02335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5559" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[112];
  assign _02337_ = _02336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5560" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[113];
  assign _02338_ = _02337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5560" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[114];
  assign _02339_ = _02338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5561" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[115];
  assign _02340_ = _02339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5561" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[116];
  assign _02341_ = _02340_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5562" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[117];
  assign _02342_ = _02341_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5562" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[118];
  assign _02343_ = _02342_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5563" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[119];
  assign _02344_ = _02343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5563" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[120];
  assign _02345_ = _02344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5564" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[121];
  assign _02346_ = _02345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5564" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[122];
  assign _02347_ = _02346_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5565" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[123];
  assign _02348_ = _02347_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5565" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[124];
  assign _02349_ = _02348_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5566" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[125];
  assign _02350_ = _02349_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5566" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[126];
  assign _02351_ = _02350_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5567" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[127];
  assign _02352_ = _02351_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5567" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[128];
  assign _02353_ = _02352_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5568" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[129];
  assign _02354_ = _02353_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5568" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[130];
  assign _02355_ = _02354_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5569" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[131];
  assign _02356_ = _02355_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5569" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[132];
  assign _02357_ = _02356_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5570" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[133];
  assign _02358_ = _02357_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5570" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[134];
  assign _02359_ = _02358_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5571" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[135];
  assign _02360_ = _02359_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5571" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[136];
  assign _02361_ = _02360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5572" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[137];
  assign _02362_ = _02361_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5572" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[138];
  assign _02363_ = _02362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5573" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[139];
  assign _02364_ = _02363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5573" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[140];
  assign _02365_ = _02364_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5574" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[141];
  assign _02366_ = _02365_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5574" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[142];
  assign _02367_ = _02366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5575" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[143];
  assign _02368_ = _02367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5575" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[144];
  assign _02369_ = _02368_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5576" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[145];
  assign _02370_ = _02369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5576" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[146];
  assign _02371_ = _02370_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5577" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[147];
  assign _02372_ = _02371_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5577" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[148];
  assign _02373_ = _02372_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5578" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[149];
  assign _02374_ = _02373_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5578" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[150];
  assign _02375_ = _02374_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5579" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[151];
  assign _02376_ = _02375_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5579" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[152];
  assign _02377_ = _02376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5580" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[153];
  assign _02378_ = _02377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5580" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[154];
  assign _02379_ = _02378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5581" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[155];
  assign _02380_ = _02379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5581" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[156];
  assign _02381_ = _02380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5582" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[157];
  assign _02382_ = _02381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5582" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[158];
  assign _02383_ = _02382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5583" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[159];
  assign _02384_ = _02383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5583" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[160];
  assign _02385_ = _02384_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5584" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[161];
  assign _02386_ = _02385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5584" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[162];
  assign _02387_ = _02386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5585" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[163];
  assign _02388_ = _02387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5585" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[164];
  assign _02389_ = _02388_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5586" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[165];
  assign _02390_ = _02389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5586" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[166];
  assign _02391_ = _02390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5587" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[167];
  assign _02392_ = _02391_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5587" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[168];
  assign _02393_ = _02392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5588" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[169];
  assign _02394_ = _02393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5588" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[170];
  assign _02395_ = _02394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5589" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[171];
  assign _02396_ = _02395_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5589" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[172];
  assign _02397_ = _02396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5590" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[173];
  assign _02398_ = _02397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5590" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[174];
  assign _02399_ = _02398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5591" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[175];
  assign _02400_ = _02399_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5591" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[176];
  assign _02401_ = _02400_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5592" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[177];
  assign _02402_ = _02401_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5592" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[178];
  assign _02403_ = _02402_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5593" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[179];
  assign _02404_ = _02403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5593" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[180];
  assign _02405_ = _02404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5594" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[181];
  assign _02406_ = _02405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5594" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[182];
  assign _02407_ = _02406_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5595" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[183];
  assign _02408_ = _02407_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5595" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[184];
  assign _02409_ = _02408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5596" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[185];
  assign _02410_ = _02409_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5596" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[186];
  assign _02411_ = _02410_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5597" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[187];
  assign _02412_ = _02411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5597" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[188];
  assign _02413_ = _02412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5598" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[189];
  assign _02414_ = _02413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5598" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[190];
  assign _02415_ = _02414_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5599" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[191];
  assign _02416_ = _02415_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5599" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[192];
  assign _02417_ = _02416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5600" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[193];
  assign _02418_ = _02417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5600" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[194];
  assign _02419_ = _02418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5601" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[195];
  assign _02420_ = _02419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5601" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[196];
  assign _02421_ = _02420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5602" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[197];
  assign _02422_ = _02421_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5602" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[198];
  assign _02423_ = _02422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5603" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[199];
  assign _02424_ = _02423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5603" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[200];
  assign _02425_ = _02424_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5604" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[201];
  assign _02426_ = _02425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5604" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[202];
  assign _02427_ = _02426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5605" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[203];
  assign _02428_ = _02427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5605" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[204];
  assign _02429_ = _02428_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5606" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[205];
  assign _02430_ = _02429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5606" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[206];
  assign _02431_ = _02430_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5607" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[207];
  assign _02432_ = _02431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5607" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[208];
  assign _02433_ = _02432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5608" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[209];
  assign _02434_ = _02433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5608" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[210];
  assign _02435_ = _02434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5609" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[211];
  assign _02436_ = _02435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5609" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[212];
  assign _02437_ = _02436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5610" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[213];
  assign _02438_ = _02437_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5610" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[214];
  assign _02439_ = _02438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5611" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[215];
  assign _02440_ = _02439_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5611" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[216];
  assign _02441_ = _02440_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5612" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[217];
  assign _02442_ = _02441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5612" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[218];
  assign _02443_ = _02442_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5613" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[219];
  assign _02444_ = _02443_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5613" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[220];
  assign _02445_ = _02444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5614" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[221];
  assign _02446_ = _02445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5614" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[222];
  assign _02447_ = _02446_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5615" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[223];
  assign _02448_ = _02447_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5615" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[224];
  assign _02449_ = _02448_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5616" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[225];
  assign _02450_ = _02449_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5616" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[226];
  assign _02451_ = _02450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5617" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[227];
  assign _02452_ = _02451_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5617" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[228];
  assign _02453_ = _02452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5618" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[229];
  assign _02454_ = _02453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5618" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[230];
  assign _02455_ = _02454_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5619" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[231];
  assign _02456_ = _02455_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5619" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[232];
  assign _02457_ = _02456_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5620" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[233];
  assign _02458_ = _02457_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5620" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[234];
  assign _02459_ = _02458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5621" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[235];
  assign _02460_ = _02459_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5621" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[236];
  assign _02461_ = _02460_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5622" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[237];
  assign _02462_ = _02461_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5622" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[238];
  assign _02463_ = _02462_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5623" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[239];
  assign _02464_ = _02463_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5623" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[240];
  assign _02465_ = _02464_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5624" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[241];
  assign _02466_ = _02465_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5624" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[242];
  assign _02467_ = _02466_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5625" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[243];
  assign _02468_ = _02467_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5625" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[244];
  assign _02469_ = _02468_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5626" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[245];
  assign _02470_ = _02469_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5626" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[246];
  assign _02471_ = _02470_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5627" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[247];
  assign _02472_ = _02471_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5627" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[248];
  assign _02473_ = _02472_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5628" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[249];
  assign _02474_ = _02473_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5628" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[250];
  assign _02475_ = _02474_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5629" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[251];
  assign _02476_ = _02475_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5629" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[252];
  assign _02477_ = _02476_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5630" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[253];
  assign _02478_ = _02477_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5630" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[254];
  assign _02479_ = _02478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5631" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[255];
  assign _02480_ = _02479_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5631" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[256];
  assign _02481_ = _02480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5632" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[257];
  assign _02482_ = _02481_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5632" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[258];
  assign _02483_ = _02482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5633" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[259];
  assign _02484_ = _02483_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5633" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[260];
  assign _02485_ = _02484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5634" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[261];
  assign _02486_ = _02485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5634" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[262];
  assign _02487_ = _02486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5635" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[263];
  assign _02488_ = _02487_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5635" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[264];
  assign _02489_ = _02488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5636" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[265];
  assign _02490_ = _02489_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5636" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[266];
  assign _02491_ = _02490_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5637" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[267];
  assign _02492_ = _02491_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5637" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[268];
  assign _02493_ = _02492_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5638" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[269];
  assign _02494_ = _02493_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5638" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[270];
  assign _02495_ = _02494_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5639" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[271];
  assign _02496_ = _02495_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5639" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[272];
  assign _02497_ = _02496_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5640" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[273];
  assign _02498_ = _02497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5640" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[274];
  assign _02499_ = _02498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5641" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[275];
  assign _02500_ = _02499_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5641" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[276];
  assign _02501_ = _02500_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5642" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[277];
  assign _02502_ = _02501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5642" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[278];
  assign _02503_ = _02502_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5643" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[279];
  assign _02504_ = _02503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5643" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[280];
  assign _02505_ = _02504_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5644" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[281];
  assign _02506_ = _02505_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5644" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[282];
  assign _02507_ = _02506_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5645" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[283];
  assign _02508_ = _02507_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5645" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[284];
  assign _02509_ = _02508_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5646" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[285];
  assign _02510_ = _02509_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5646" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[286];
  assign _02511_ = _02510_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5647" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[287];
  assign _02512_ = _02511_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5647" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[288];
  assign _02513_ = _02512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5648" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[289];
  assign _02514_ = _02513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5648" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[290];
  assign _02515_ = _02514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5649" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[291];
  assign _02516_ = _02515_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5649" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[292];
  assign _02517_ = _02516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5650" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[293];
  assign _02518_ = _02517_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5650" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[294];
  assign _02519_ = _02518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5651" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[295];
  assign _02520_ = _02519_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5651" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[296];
  assign _02521_ = _02520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5652" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[297];
  assign _02522_ = _02521_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5652" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[298];
  assign _02523_ = _02522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5653" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[299];
  assign _02524_ = _02523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5653" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[300];
  assign _02525_ = _02524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5654" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[301];
  assign _02526_ = _02525_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5654" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[302];
  assign _02527_ = _02526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5655" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[303];
  assign _02528_ = _02527_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5655" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[304];
  assign _02529_ = _02528_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5656" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[305];
  assign _02530_ = _02529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5656" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[306];
  assign _02531_ = _02530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5657" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[307];
  assign _02532_ = _02531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5657" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[308];
  assign _02533_ = _02532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5658" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[309];
  assign _02534_ = _02533_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5658" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[310];
  assign _02535_ = _02534_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5659" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[311];
  assign _02536_ = _02535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5659" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[312];
  assign _02537_ = _02536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5660" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[313];
  assign _02538_ = _02537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5660" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[314];
  assign _02539_ = _02538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5661" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[315];
  assign _02540_ = _02539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5661" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[316];
  assign _02541_ = _02540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5662" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[317];
  assign _02542_ = _02541_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5662" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[318];
  assign _02543_ = _02542_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5663" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[319];
  assign _02544_ = _02543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5663" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[320];
  assign _02545_ = _02544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5664" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[321];
  assign _02546_ = _02545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5664" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[322];
  assign _02547_ = _02546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5665" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[323];
  assign _02548_ = _02547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5665" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[324];
  assign _02549_ = _02548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5666" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[325];
  assign _02550_ = _02549_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5666" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[326];
  assign _02551_ = _02550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5667" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[327];
  assign _02552_ = _02551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5667" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[328];
  assign _02553_ = _02552_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5668" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[329];
  assign _02554_ = _02553_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5668" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[330];
  assign _02555_ = _02554_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5669" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[331];
  assign _02556_ = _02555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5669" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[332];
  assign _02557_ = _02556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5670" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[333];
  assign _02558_ = _02557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5670" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[334];
  assign _02559_ = _02558_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5671" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[335];
  assign _02560_ = _02559_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5671" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[336];
  assign _02561_ = _02560_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5672" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[337];
  assign _02562_ = _02561_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5672" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[338];
  assign _02563_ = _02562_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5673" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[339];
  assign _02564_ = _02563_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5673" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[340];
  assign _02565_ = _02564_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5674" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[341];
  assign _02566_ = _02565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5674" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[342];
  assign _02567_ = _02566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5675" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[343];
  assign _02568_ = _02567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5675" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[344];
  assign _02569_ = _02568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5676" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[345];
  assign _02570_ = _02569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5676" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[346];
  assign _02571_ = _02570_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5677" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[347];
  assign _02572_ = _02571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5677" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[348];
  assign _02573_ = _02572_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5678" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[349];
  assign _02574_ = _02573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5678" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[350];
  assign _02575_ = _02574_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5679" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[351];
  assign _02576_ = _02575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5679" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[352];
  assign _02577_ = _02576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5680" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[353];
  assign _02578_ = _02577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5680" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[354];
  assign _02579_ = _02578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5681" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[355];
  assign _02580_ = _02579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5681" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[356];
  assign _02581_ = _02580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5682" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[357];
  assign _02582_ = _02581_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5682" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[358];
  assign _02583_ = _02582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5683" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[359];
  assign _02584_ = _02583_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5683" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[360];
  assign _02585_ = _02584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5684" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[361];
  assign _02586_ = _02585_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5684" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[362];
  assign _02587_ = _02586_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5685" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[363];
  assign _02588_ = _02587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5685" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[364];
  assign _02589_ = _02588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5686" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[365];
  assign _02590_ = _02589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5686" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[366];
  assign _02591_ = _02590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5687" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[367];
  assign _02592_ = _02591_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5687" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[368];
  assign _02593_ = _02592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5688" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[369];
  assign _02594_ = _02593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5688" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[370];
  assign _02595_ = _02594_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5689" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[371];
  assign _02596_ = _02595_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5689" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[372];
  assign _02597_ = _02596_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5690" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[373];
  assign _02598_ = _02597_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5690" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[374];
  assign _02599_ = _02598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5691" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[375];
  assign _02600_ = _02599_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5691" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[376];
  assign _02601_ = _02600_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5692" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[377];
  assign _02602_ = _02601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5692" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[378];
  assign _02603_ = _02602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5693" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[379];
  assign _02604_ = _02603_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5693" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[380];
  assign _02605_ = _02604_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5694" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[381];
  assign _02606_ = _02605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5694" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[382];
  assign _02607_ = _02606_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5695" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[383];
  assign _02608_ = _02607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5695" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[384];
  assign _02609_ = _02608_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5696" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[385];
  assign _02610_ = _02609_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5696" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[386];
  assign _02611_ = _02610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5697" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[387];
  assign _02612_ = _02611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5697" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[388];
  assign _02613_ = _02612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5698" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[389];
  assign _02614_ = _02613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5698" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[390];
  assign _02615_ = _02614_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5699" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[391];
  assign _02616_ = _02615_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5699" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[392];
  assign _02617_ = _02616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5700" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[393];
  assign _02618_ = _02617_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5700" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[394];
  assign _02619_ = _02618_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5701" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[395];
  assign _02620_ = _02619_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5701" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[396];
  assign _02621_ = _02620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5702" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[397];
  assign _02622_ = _02621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5702" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[398];
  assign _02623_ = _02622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5703" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[399];
  assign _02624_ = _02623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5703" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[400];
  assign _02625_ = _02624_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5704" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[401];
  assign _02626_ = _02625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5704" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[402];
  assign _02627_ = _02626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5705" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[403];
  assign _02628_ = _02627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5705" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[404];
  assign _02629_ = _02628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5706" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[405];
  assign _02630_ = _02629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5706" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[406];
  assign _02631_ = _02630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5707" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[407];
  assign _02632_ = _02631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5707" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[408];
  assign _02633_ = _02632_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5708" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[409];
  assign _02634_ = _02633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5708" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[410];
  assign _02635_ = _02634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5709" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[411];
  assign _02636_ = _02635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5709" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[412];
  assign _02637_ = _02636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5710" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[413];
  assign _02638_ = _02637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5710" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[414];
  assign _02639_ = _02638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5711" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[415];
  assign _02640_ = _02639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5711" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[416];
  assign _02641_ = _02640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5712" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[417];
  assign _02642_ = _02641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5712" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[418];
  assign _02643_ = _02642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5713" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[419];
  assign _02644_ = _02643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5713" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[420];
  assign _02645_ = _02644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5714" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[421];
  assign _02646_ = _02645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5714" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[422];
  assign _02647_ = _02646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5715" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[423];
  assign _02648_ = _02647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5715" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[424];
  assign _02649_ = _02648_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5716" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[425];
  assign _02650_ = _02649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5716" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[426];
  assign _02651_ = _02650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5717" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[427];
  assign _02652_ = _02651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5717" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[428];
  assign _02653_ = _02652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5718" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[429];
  assign _02654_ = _02653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5718" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[430];
  assign _02655_ = _02654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5719" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[431];
  assign _02656_ = _02655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5719" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[432];
  assign _02657_ = _02656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5720" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[433];
  assign _02658_ = _02657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5720" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[434];
  assign _02659_ = _02658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5721" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[435];
  assign _02660_ = _02659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5721" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[436];
  assign _02661_ = _02660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5722" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[437];
  assign _02662_ = _02661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5722" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[438];
  assign _02663_ = _02662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5723" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[439];
  assign _02664_ = _02663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5723" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[440];
  assign _02665_ = _02664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5724" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[441];
  assign _02666_ = _02665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5724" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[442];
  assign _02667_ = _02666_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5725" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[443];
  assign _02668_ = _02667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5725" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[444];
  assign _02669_ = _02668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5726" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[445];
  assign _02670_ = _02669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5726" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[446];
  assign _02671_ = _02670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5727" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[447];
  assign _02672_ = _02671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5727" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[448];
  assign _02673_ = _02672_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5728" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[449];
  assign _02674_ = _02673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5728" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[450];
  assign _02675_ = _02674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5729" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[451];
  assign _02676_ = _02675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5729" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[452];
  assign _02677_ = _02676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5730" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[453];
  assign _02678_ = _02677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5730" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[454];
  assign _02679_ = _02678_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5731" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[455];
  assign _02680_ = _02679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5731" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[456];
  assign _02681_ = _02680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5732" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[457];
  assign _02682_ = _02681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5732" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[458];
  assign _02683_ = _02682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5733" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[459];
  assign _02684_ = _02683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5733" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[460];
  assign _02685_ = _02684_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5734" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[461];
  assign _02686_ = _02685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5734" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[462];
  assign _02687_ = _02686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5735" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[463];
  assign _02688_ = _02687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5735" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[464];
  assign _02689_ = _02688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5736" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[465];
  assign _02690_ = _02689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5736" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[466];
  assign _02691_ = _02690_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5737" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[467];
  assign _02692_ = _02691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5737" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[468];
  assign _02693_ = _02692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5738" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[469];
  assign _02694_ = _02693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5738" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[470];
  assign _02695_ = _02694_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5739" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[471];
  assign _02696_ = _02695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5739" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[472];
  assign _02697_ = _02696_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5740" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[473];
  assign _02698_ = _02697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5740" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[474];
  assign _02699_ = _02698_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5741" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[475];
  assign _02700_ = _02699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5741" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[476];
  assign _02701_ = _02700_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5742" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[477];
  assign _02702_ = _02701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5742" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[478];
  assign _02703_ = _02702_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5743" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[479];
  assign _02704_ = _02703_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5743" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[480];
  assign _02705_ = _02704_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5744" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[481];
  assign _02706_ = _02705_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5744" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[482];
  assign _02707_ = _02706_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5745" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[483];
  assign _02708_ = _02707_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5745" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[484];
  assign _02709_ = _02708_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5746" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[485];
  assign _02710_ = _02709_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5746" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[486];
  assign _02711_ = _02710_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5747" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[487];
  assign _02712_ = _02711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5747" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[488];
  assign _02713_ = _02712_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5748" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[489];
  assign _02714_ = _02713_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5748" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[490];
  assign _02715_ = _02714_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5749" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[491];
  assign _02716_ = _02715_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5749" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[492];
  assign _02717_ = _02716_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5750" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[493];
  assign _02718_ = _02717_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5750" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[494];
  assign _02719_ = _02718_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5751" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[495];
  assign _02720_ = _02719_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5751" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[496];
  assign _02721_ = _02720_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5752" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[497];
  assign _02722_ = _02721_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5752" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[498];
  assign _02723_ = _02722_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5753" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[499];
  assign _02724_ = _02723_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5753" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[500];
  assign _02725_ = _02724_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5754" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[501];
  assign _02726_ = _02725_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5754" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[502];
  assign _02727_ = _02726_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5755" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[503];
  assign _02728_ = _02727_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5755" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[504];
  assign _02729_ = _02728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5756" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[505];
  assign _02730_ = _02729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5756" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[506];
  assign _02731_ = _02730_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5757" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[507];
  assign _02732_ = _02731_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5757" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[508];
  assign _02733_ = _02732_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5758" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[509];
  assign _02734_ = _02733_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5758" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[510];
  assign _02735_ = _02734_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5759" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[511];
  assign _02736_ = _02735_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5759" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[512];
  assign _02737_ = _02736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5760" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[513];
  assign _02738_ = _02737_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5760" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[514];
  assign _02739_ = _02738_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5761" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[515];
  assign _02740_ = _02739_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5761" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[516];
  assign _02741_ = _02740_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5762" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[517];
  assign _02742_ = _02741_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5762" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[518];
  assign _02743_ = _02742_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5763" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[519];
  assign _02744_ = _02743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5763" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[520];
  assign _02745_ = _02744_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5764" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[521];
  assign _02746_ = _02745_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5764" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[522];
  assign _02747_ = _02746_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5765" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[523];
  assign _02748_ = _02747_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5765" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[524];
  assign _02749_ = _02748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5766" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[525];
  assign _02750_ = _02749_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5766" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[526];
  assign _02751_ = _02750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5767" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[527];
  assign _02752_ = _02751_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5767" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[528];
  assign _02753_ = _02752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5768" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[529];
  assign _02754_ = _02753_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5768" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[530];
  assign _02755_ = _02754_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5769" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[531];
  assign _02756_ = _02755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5769" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[532];
  assign _02757_ = _02756_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5770" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[533];
  assign _02758_ = _02757_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5770" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[534];
  assign _02759_ = _02758_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5771" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[535];
  assign _02760_ = _02759_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5771" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[536];
  assign _02761_ = _02760_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5772" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[537];
  assign _02762_ = _02761_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5772" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[538];
  assign _02763_ = _02762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5773" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[539];
  assign _02764_ = _02763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5773" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[540];
  assign _02765_ = _02764_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5774" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[541];
  assign _02766_ = _02765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5774" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[542];
  assign _02767_ = _02766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5775" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[543];
  assign _02768_ = _02767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5775" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[544];
  assign _02769_ = _02768_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5776" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[545];
  assign _02770_ = _02769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5776" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[546];
  assign _02771_ = _02770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5777" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[547];
  assign _02772_ = _02771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5777" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[548];
  assign _02773_ = _02772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5778" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[549];
  assign _02774_ = _02773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5778" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[550];
  assign _02775_ = _02774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5779" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[551];
  assign _02776_ = _02775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5779" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[552];
  assign _02777_ = _02776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5780" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[553];
  assign _02778_ = _02777_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5780" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[554];
  assign _02779_ = _02778_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5781" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[555];
  assign _02780_ = _02779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5781" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[556];
  assign _02781_ = _02780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5782" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[557];
  assign _02782_ = _02781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5782" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[558];
  assign _02783_ = _02782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5783" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[559];
  assign _02784_ = _02783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5783" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[560];
  assign _02785_ = _02784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5784" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[561];
  assign _02786_ = _02785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5784" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[562];
  assign _02787_ = _02786_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5785" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[563];
  assign _02788_ = _02787_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5785" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[564];
  assign _02789_ = _02788_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5786" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[565];
  assign _02790_ = _02789_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5786" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[566];
  assign _02791_ = _02790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5787" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[567];
  assign _02792_ = _02791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5787" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[568];
  assign _02793_ = _02792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5788" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[569];
  assign _02794_ = _02793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5788" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[570];
  assign _02795_ = _02794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5789" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[571];
  assign _02796_ = _02795_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5789" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[572];
  assign _02797_ = _02796_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5790" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[573];
  assign _02798_ = _02797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5790" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[574];
  assign _02799_ = _02798_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5791" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[575];
  assign _02800_ = _02799_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5791" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[576];
  assign _02801_ = _02800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5792" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[577];
  assign _02802_ = _02801_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5792" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[578];
  assign _02803_ = _02802_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5793" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[579];
  assign _02804_ = _02803_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5793" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[580];
  assign _02805_ = _02804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5794" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[581];
  assign _02806_ = _02805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5794" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[582];
  assign _02807_ = _02806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5795" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[583];
  assign _02808_ = _02807_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5795" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[584];
  assign _02809_ = _02808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5796" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[585];
  assign _02810_ = _02809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5796" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[586];
  assign _02811_ = _02810_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5797" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[587];
  assign _02812_ = _02811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5797" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[588];
  assign _02813_ = _02812_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5798" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[589];
  assign _02814_ = _02813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5798" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[590];
  assign _02815_ = _02814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5799" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[591];
  assign _02816_ = _02815_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5799" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[592];
  assign _02817_ = _02816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5800" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[593];
  assign _02818_ = _02817_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5800" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[594];
  assign _02819_ = _02818_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5801" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[595];
  assign _02820_ = _02819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5801" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[596];
  assign _02821_ = _02820_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5802" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[597];
  assign _02822_ = _02821_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5802" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[598];
  assign _02823_ = _02822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5803" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[599];
  assign _02824_ = _02823_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5803" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[600];
  assign _02825_ = _02824_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5804" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[601];
  assign _02826_ = _02825_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5804" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[602];
  assign _02827_ = _02826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5805" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[603];
  assign _02828_ = _02827_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5805" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[604];
  assign _02829_ = _02828_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5806" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[605];
  assign _02830_ = _02829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5806" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[606];
  assign _02831_ = _02830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5807" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[607];
  assign _02832_ = _02831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5807" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[608];
  assign _02833_ = _02832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5808" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[609];
  assign _02834_ = _02833_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5808" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[610];
  assign _02835_ = _02834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5809" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[611];
  assign _02836_ = _02835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5809" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[612];
  assign _02837_ = _02836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5810" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[613];
  assign _02838_ = _02837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5810" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[614];
  assign _02839_ = _02838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5811" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[615];
  assign _02840_ = _02839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5811" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[616];
  assign _02841_ = _02840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5812" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[617];
  assign _02842_ = _02841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5812" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[618];
  assign _02843_ = _02842_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5813" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[619];
  assign _02844_ = _02843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5813" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[620];
  assign _02845_ = _02844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5814" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[621];
  assign _02846_ = _02845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5814" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[622];
  assign _02847_ = _02846_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5815" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[623];
  assign _02848_ = _02847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5815" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[624];
  assign _02849_ = _02848_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5816" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[625];
  assign _02850_ = _02849_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5816" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[626];
  assign _02851_ = _02850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5817" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[627];
  assign _02852_ = _02851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5817" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[628];
  assign _02853_ = _02852_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5818" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[629];
  assign _02854_ = _02853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5818" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[630];
  assign _02855_ = _02854_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5819" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[631];
  assign _02856_ = _02855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5819" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[632];
  assign _02857_ = _02856_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5820" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[633];
  assign _02858_ = _02857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5820" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[634];
  assign _02859_ = _02858_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5821" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[635];
  assign _02860_ = _02859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5821" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[636];
  assign _02861_ = _02860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5822" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[637];
  assign _02862_ = _02861_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5822" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[638];
  assign _02863_ = _02862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5823" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[639];
  assign _02864_ = _02863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5823" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[640];
  assign _02865_ = _02864_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5824" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[641];
  assign _02866_ = _02865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5824" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[642];
  assign _02867_ = _02866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5825" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[643];
  assign _02868_ = _02867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5825" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[644];
  assign _02869_ = _02868_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5826" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[645];
  assign _02870_ = _02869_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5826" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[646];
  assign _02871_ = _02870_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5827" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[647];
  assign _02872_ = _02871_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5827" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[648];
  assign _02873_ = _02872_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5828" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[649];
  assign _02874_ = _02873_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5828" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[650];
  assign _02875_ = _02874_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5829" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[651];
  assign _02876_ = _02875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5829" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[652];
  assign _02877_ = _02876_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5830" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[653];
  assign _02878_ = _02877_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5830" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[654];
  assign _02879_ = _02878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5831" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[655];
  assign _02880_ = _02879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5831" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[656];
  assign _02881_ = _02880_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5832" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[657];
  assign _02882_ = _02881_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5832" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[658];
  assign _02883_ = _02882_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5833" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[659];
  assign _02884_ = _02883_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5833" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[660];
  assign _02885_ = _02884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5834" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[661];
  assign _02886_ = _02885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5834" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[662];
  assign _02887_ = _02886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5835" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[663];
  assign _02888_ = _02887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5835" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[664];
  assign _02889_ = _02888_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5836" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[665];
  assign _02890_ = _02889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5836" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[666];
  assign _02891_ = _02890_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5837" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[667];
  assign _02892_ = _02891_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5837" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[668];
  assign _02893_ = _02892_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5838" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[669];
  assign _02894_ = _02893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5838" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[670];
  assign _02895_ = _02894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5839" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[671];
  assign _02896_ = _02895_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5839" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[672];
  assign _02897_ = _02896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5840" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[673];
  assign _02898_ = _02897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5840" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[674];
  assign _02899_ = _02898_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5841" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[675];
  assign _02900_ = _02899_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5841" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[676];
  assign _02901_ = _02900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5842" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[677];
  assign _02902_ = _02901_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5842" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[678];
  assign _02903_ = _02902_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5843" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[679];
  assign _02904_ = _02903_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5843" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[680];
  assign _02905_ = _02904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5844" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[681];
  assign _02906_ = _02905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5844" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[682];
  assign _02907_ = _02906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5845" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[683];
  assign _02908_ = _02907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5845" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[684];
  assign _02909_ = _02908_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5846" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[685];
  assign _02910_ = _02909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5846" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[686];
  assign _02911_ = _02910_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5847" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[687];
  assign _02912_ = _02911_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5847" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[688];
  assign _02913_ = _02912_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5848" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[689];
  assign _02914_ = _02913_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5848" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[690];
  assign _02915_ = _02914_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5849" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[691];
  assign _02916_ = _02915_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5849" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[692];
  assign _02917_ = _02916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5850" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[693];
  assign _02918_ = _02917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5850" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[694];
  assign _02919_ = _02918_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5851" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[695];
  assign _02920_ = _02919_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5851" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[696];
  assign _02921_ = _02920_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5852" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[697];
  assign _02922_ = _02921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5852" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[698];
  assign _02923_ = _02922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5853" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[699];
  assign _02924_ = _02923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5853" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[700];
  assign _02925_ = _02924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5854" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[701];
  assign _02926_ = _02925_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5854" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[702];
  assign _02927_ = _02926_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5855" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[703];
  assign _02928_ = _02927_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5855" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[704];
  assign _02929_ = _02928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5856" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[705];
  assign _02930_ = _02929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5856" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[706];
  assign _02931_ = _02930_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5857" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[707];
  assign _02932_ = _02931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5857" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[708];
  assign _02933_ = _02932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5858" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[709];
  assign _02934_ = _02933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5858" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[710];
  assign _02935_ = _02934_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5859" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[711];
  assign _02936_ = _02935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5859" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[712];
  assign _02937_ = _02936_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5860" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[713];
  assign _02938_ = _02937_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5860" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[714];
  assign _02939_ = _02938_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5861" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[715];
  assign _02940_ = _02939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5861" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[716];
  assign _02941_ = _02940_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5862" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[717];
  assign _02942_ = _02941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5862" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[718];
  assign _02943_ = _02942_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5863" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[719];
  assign _02944_ = _02943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5863" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[720];
  assign _02945_ = _02944_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5864" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[721];
  assign _02946_ = _02945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5864" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[722];
  assign _02947_ = _02946_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5865" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[723];
  assign _02948_ = _02947_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5865" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[724];
  assign _02949_ = _02948_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5866" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[725];
  assign _02950_ = _02949_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5866" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[726];
  assign _02951_ = _02950_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5867" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[727];
  assign _02952_ = _02951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5867" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[728];
  assign _02953_ = _02952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5868" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[729];
  assign _02954_ = _02953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5868" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[730];
  assign _02955_ = _02954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5869" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[731];
  assign _02956_ = _02955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5869" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[732];
  assign _02957_ = _02956_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5870" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[733];
  assign _02958_ = _02957_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5870" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[734];
  assign _02959_ = _02958_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5871" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[735];
  assign _02960_ = _02959_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5871" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[736];
  assign _02961_ = _02960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5872" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[737];
  assign _02962_ = _02961_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5872" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[738];
  assign _02963_ = _02962_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5873" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[739];
  assign _02964_ = _02963_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5873" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[740];
  assign _02965_ = _02964_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5874" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[741];
  assign _02966_ = _02965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5874" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[742];
  assign _02967_ = _02966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5875" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[743];
  assign _02968_ = _02967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5875" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[744];
  assign _02969_ = _02968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5876" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[745];
  assign _02970_ = _02969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5876" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[746];
  assign _02971_ = _02970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5877" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[747];
  assign _02972_ = _02971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5877" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[748];
  assign _02973_ = _02972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5878" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[749];
  assign _02974_ = _02973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5878" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[750];
  assign _02975_ = _02974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5879" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[751];
  assign _02976_ = _02975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5879" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[752];
  assign _02977_ = _02976_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5880" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[753];
  assign _02978_ = _02977_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5880" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[754];
  assign _02979_ = _02978_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5881" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[755];
  assign _02980_ = _02979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5881" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[756];
  assign _02981_ = _02980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5882" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[757];
  assign _02982_ = _02981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5882" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[758];
  assign _02983_ = _02982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5883" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[759];
  assign _02984_ = _02983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5883" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[760];
  assign _02985_ = _02984_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5884" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[761];
  assign _02986_ = _02985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5884" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[762];
  assign _02987_ = _02986_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5885" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[763];
  assign _02988_ = _02987_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5885" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[764];
  assign _02989_ = _02988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5886" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[765];
  assign _02990_ = _02989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5886" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[766];
  assign _02991_ = _02990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5887" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[767];
  assign _02992_ = _02991_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5887" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[768];
  assign _02993_ = _02992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5888" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[769];
  assign _02994_ = _02993_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5888" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[770];
  assign _02995_ = _02994_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5889" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[771];
  assign _02996_ = _02995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5889" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[772];
  assign _02997_ = _02996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5890" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[773];
  assign _02998_ = _02997_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5890" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[774];
  assign _02999_ = _02998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5891" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[775];
  assign _03000_ = _02999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5891" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[776];
  assign _03001_ = _03000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5892" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[777];
  assign _03002_ = _03001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5892" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[778];
  assign _03003_ = _03002_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5893" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[779];
  assign _03004_ = _03003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5893" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[780];
  assign _03005_ = _03004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5894" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[781];
  assign _03006_ = _03005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5894" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[782];
  assign _03007_ = _03006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5895" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[783];
  assign _03008_ = _03007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5895" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[784];
  assign _03009_ = _03008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5896" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[785];
  assign _03010_ = _03009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5896" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[786];
  assign _03011_ = _03010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5897" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[787];
  assign _03012_ = _03011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5897" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[788];
  assign _03013_ = _03012_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5898" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[789];
  assign _03014_ = _03013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5898" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[790];
  assign _03015_ = _03014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5899" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[791];
  assign _03016_ = _03015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5899" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[792];
  assign _03017_ = _03016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5900" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[793];
  assign _03018_ = _03017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5900" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[794];
  assign _03019_ = _03018_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5901" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[795];
  assign _03020_ = _03019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5901" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[796];
  assign _03021_ = _03020_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5902" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[797];
  assign _03022_ = _03021_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5902" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[798];
  assign _03023_ = _03022_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5903" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[799];
  assign _03024_ = _03023_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5903" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[800];
  assign _03025_ = _03024_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5904" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[801];
  assign _03026_ = _03025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5904" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[802];
  assign _03027_ = _03026_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5905" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[803];
  assign _03028_ = _03027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5905" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[804];
  assign _03029_ = _03028_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5906" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[805];
  assign _03030_ = _03029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5906" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[806];
  assign _03031_ = _03030_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5907" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[807];
  assign _03032_ = _03031_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5907" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[808];
  assign _03033_ = _03032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5908" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[809];
  assign _03034_ = _03033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5908" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[810];
  assign _03035_ = _03034_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5909" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[811];
  assign _03036_ = _03035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5909" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[812];
  assign _03037_ = _03036_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5910" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[813];
  assign _03038_ = _03037_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5910" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[814];
  assign _03039_ = _03038_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5911" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[815];
  assign _03040_ = _03039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5911" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[816];
  assign _03041_ = _03040_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5912" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[817];
  assign _03042_ = _03041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5912" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[818];
  assign _03043_ = _03042_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5913" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[819];
  assign _03044_ = _03043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5913" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[820];
  assign _03045_ = _03044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5914" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[821];
  assign _03046_ = _03045_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5914" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[822];
  assign _03047_ = _03046_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5915" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[823];
  assign _03048_ = _03047_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5915" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[824];
  assign _03049_ = _03048_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5916" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[825];
  assign _03050_ = _03049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5916" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[826];
  assign _03051_ = _03050_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5917" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[827];
  assign _03052_ = _03051_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5917" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[828];
  assign _03053_ = _03052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5918" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[829];
  assign _03054_ = _03053_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5918" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[830];
  assign _03055_ = _03054_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5919" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[831];
  assign _03056_ = _03055_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5919" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[832];
  assign _03057_ = _03056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5920" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[833];
  assign _03058_ = _03057_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5920" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[834];
  assign _03059_ = _03058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5921" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[835];
  assign _03060_ = _03059_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5921" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[836];
  assign _03061_ = _03060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5922" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[837];
  assign _03062_ = _03061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5922" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[838];
  assign _03063_ = _03062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5923" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[839];
  assign _03064_ = _03063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5923" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[840];
  assign _03065_ = _03064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5924" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[841];
  assign _03066_ = _03065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5924" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[842];
  assign _03067_ = _03066_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5925" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[843];
  assign _03068_ = _03067_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5925" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[844];
  assign _03069_ = _03068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5926" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[845];
  assign _03070_ = _03069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5926" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[846];
  assign _03071_ = _03070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5927" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[847];
  assign _03072_ = _03071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5927" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[848];
  assign _03073_ = _03072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5928" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[849];
  assign _03074_ = _03073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5928" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[850];
  assign _03075_ = _03074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5929" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[851];
  assign _03076_ = _03075_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5929" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[852];
  assign _03077_ = _03076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5930" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[853];
  assign _03078_ = _03077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5930" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[854];
  assign _03079_ = _03078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5931" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[855];
  assign _03080_ = _03079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5931" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[856];
  assign _03081_ = _03080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5932" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[857];
  assign _03082_ = _03081_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5932" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[858];
  assign _03083_ = _03082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5933" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[859];
  assign _03084_ = _03083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5933" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[860];
  assign _03085_ = _03084_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5934" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[861];
  assign _03086_ = _03085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5934" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[862];
  assign _03087_ = _03086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5935" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[863];
  assign _03088_ = _03087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5935" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[864];
  assign _03089_ = _03088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5936" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[865];
  assign _03090_ = _03089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5936" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[866];
  assign _03091_ = _03090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5937" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[867];
  assign _03092_ = _03091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5937" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[868];
  assign _03093_ = _03092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5938" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[869];
  assign _03094_ = _03093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5938" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[870];
  assign _03095_ = _03094_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5939" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[871];
  assign _03096_ = _03095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5939" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[872];
  assign _03097_ = _03096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5940" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[873];
  assign _03098_ = _03097_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5940" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[874];
  assign _03099_ = _03098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5941" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[875];
  assign _03100_ = _03099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5941" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[876];
  assign _03101_ = _03100_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5942" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[877];
  assign _03102_ = _03101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5942" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[878];
  assign _03103_ = _03102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5943" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[879];
  assign _03104_ = _03103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5943" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[880];
  assign _03105_ = _03104_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5944" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[881];
  assign _03106_ = _03105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5944" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[882];
  assign _03107_ = _03106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5945" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[883];
  assign _03108_ = _03107_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5945" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[884];
  assign _03109_ = _03108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5946" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[885];
  assign _03110_ = _03109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5946" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[886];
  assign _03111_ = _03110_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5947" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[887];
  assign _03112_ = _03111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5947" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[888];
  assign _03113_ = _03112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5948" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[889];
  assign _03114_ = _03113_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5948" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[890];
  assign _03115_ = _03114_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5949" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[891];
  assign _03116_ = _03115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5949" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[892];
  assign _03117_ = _03116_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5950" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[893];
  assign _03118_ = _03117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5950" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[894];
  assign _03119_ = _03118_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5951" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[895];
  assign _03120_ = _03119_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5951" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[896];
  assign _03121_ = _03120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5952" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[897];
  assign _03122_ = _03121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5952" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[898];
  assign _03123_ = _03122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5953" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[899];
  assign _03124_ = _03123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5953" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[900];
  assign _03125_ = _03124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5954" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[901];
  assign _03126_ = _03125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5954" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[902];
  assign _03127_ = _03126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5955" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[903];
  assign _03128_ = _03127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5955" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[904];
  assign _03129_ = _03128_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5956" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[905];
  assign _03130_ = _03129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5956" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[906];
  assign _03131_ = _03130_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5957" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[907];
  assign _03132_ = _03131_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5957" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[908];
  assign _03133_ = _03132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5958" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[909];
  assign _03134_ = _03133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5958" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[910];
  assign _03135_ = _03134_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5959" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[911];
  assign _03136_ = _03135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5959" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[912];
  assign _03137_ = _03136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5960" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[913];
  assign _03138_ = _03137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5960" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[914];
  assign _03139_ = _03138_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5961" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[915];
  assign _03140_ = _03139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5961" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[916];
  assign _03141_ = _03140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5962" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[917];
  assign _03142_ = _03141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5962" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[918];
  assign _03143_ = _03142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5963" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[919];
  assign _03144_ = _03143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5963" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[920];
  assign _03145_ = _03144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5964" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[921];
  assign _03146_ = _03145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5964" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[922];
  assign _03147_ = _03146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5965" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[923];
  assign _03148_ = _03147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5965" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[924];
  assign _03149_ = _03148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5966" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[925];
  assign _03150_ = _03149_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5966" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[926];
  assign _03151_ = _03150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5967" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[927];
  assign _03152_ = _03151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5967" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[928];
  assign _03153_ = _03152_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5968" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[929];
  assign _03154_ = _03153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5968" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[930];
  assign _03155_ = _03154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5969" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[931];
  assign _03156_ = _03155_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5969" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[932];
  assign _03157_ = _03156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5970" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[933];
  assign _03158_ = _03157_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5970" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[934];
  assign _03159_ = _03158_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5971" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[935];
  assign _03160_ = _03159_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5971" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[936];
  assign _03161_ = _03160_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5972" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[937];
  assign _03162_ = _03161_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5972" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[938];
  assign _03163_ = _03162_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5973" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[939];
  assign _03164_ = _03163_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5973" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[940];
  assign _03165_ = _03164_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5974" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[941];
  assign _03166_ = _03165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5974" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[942];
  assign _03167_ = _03166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5975" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[943];
  assign _03168_ = _03167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5975" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[944];
  assign _03169_ = _03168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5976" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[945];
  assign _03170_ = _03169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5976" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[946];
  assign _03171_ = _03170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5977" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[947];
  assign _03172_ = _03171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5977" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[948];
  assign _03173_ = _03172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5978" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[949];
  assign _03174_ = _03173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5978" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[950];
  assign _03175_ = _03174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5979" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[951];
  assign _03176_ = _03175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5979" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[952];
  assign _03177_ = _03176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5980" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[953];
  assign _03178_ = _03177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5980" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[954];
  assign _03179_ = _03178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5981" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[955];
  assign _03180_ = _03179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5981" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[956];
  assign _03181_ = _03180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5982" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[957];
  assign _03182_ = _03181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5982" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[958];
  assign _03183_ = _03182_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5983" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[959];
  assign _03184_ = _03183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5983" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[960];
  assign _03185_ = _03184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5984" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[961];
  assign _03186_ = _03185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5984" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[962];
  assign _03187_ = _03186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5985" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[963];
  assign _03188_ = _03187_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5985" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[964];
  assign _03189_ = _03188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5986" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[965];
  assign _03190_ = _03189_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5986" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[966];
  assign _03191_ = _03190_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5987" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[967];
  assign _03192_ = _03191_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5987" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[968];
  assign _03193_ = _03192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5988" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[969];
  assign _03194_ = _03193_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5988" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[970];
  assign _03195_ = _03194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5989" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[971];
  assign _03196_ = _03195_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5989" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[972];
  assign _03197_ = _03196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5990" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[973];
  assign _03198_ = _03197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5990" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[974];
  assign _03199_ = _03198_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5991" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[975];
  assign _03200_ = _03199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5991" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[976];
  assign _03201_ = _03200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5992" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[977];
  assign _03202_ = _03201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5992" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[978];
  assign _03203_ = _03202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5993" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[979];
  assign _03204_ = _03203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5993" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[980];
  assign _03205_ = _03204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5994" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[981];
  assign _03206_ = _03205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5994" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[982];
  assign _03207_ = _03206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5995" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[983];
  assign _03208_ = _03207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5995" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[984];
  assign _03209_ = _03208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5996" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[985];
  assign _03210_ = _03209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5996" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[986];
  assign _03211_ = _03210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5997" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[987];
  assign _03212_ = _03211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5997" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[988];
  assign _03213_ = _03212_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5998" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[989];
  assign _03214_ = _03213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5998" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[990];
  assign _03215_ = _03214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5999" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[991];
  assign _03216_ = _03215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:5999" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[992];
  assign _03217_ = _03216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6000" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[993];
  assign _03218_ = _03217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6000" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[994];
  assign _03219_ = _03218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6001" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[995];
  assign _03220_ = _03219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6001" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[996];
  assign _03221_ = _03220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6002" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[997];
  assign _03222_ = _03221_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6002" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[998];
  assign _03223_ = _03222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6003" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[999];
  assign _03224_ = _03223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6003" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1000];
  assign _03225_ = _03224_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6004" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1001];
  assign _03226_ = _03225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6004" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1002];
  assign _03227_ = _03226_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6005" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1003];
  assign _03228_ = _03227_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6005" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1004];
  assign _03229_ = _03228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6006" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1005];
  assign _03230_ = _03229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6006" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1006];
  assign _03231_ = _03230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6007" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1007];
  assign _03232_ = _03231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6007" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1008];
  assign _03233_ = _03232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6008" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1009];
  assign _03234_ = _03233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6008" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1010];
  assign _03235_ = _03234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6009" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1011];
  assign _03236_ = _03235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6009" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1012];
  assign _03237_ = _03236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6010" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1013];
  assign _03238_ = _03237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6010" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1014];
  assign _03239_ = _03238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6011" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1015];
  assign _03240_ = _03239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6011" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1016];
  assign _03241_ = _03240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6012" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1017];
  assign _03242_ = _03241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6012" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1018];
  assign _03243_ = _03242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6013" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1019];
  assign _03244_ = _03243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6013" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1020];
  assign _03245_ = _03244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6014" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva[1021];
  assign _03246_ = _03245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6014" *) _00855_;
  assign _03247_ = IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6020" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1];
  assign _03248_ = _03247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6020" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[2];
  assign _03249_ = _03248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6021" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[3];
  assign _03250_ = _03249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6021" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[4];
  assign _03251_ = _03250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6022" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[5];
  assign _03252_ = _03251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6022" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[6];
  assign _03253_ = _03252_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6023" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[7];
  assign _03254_ = _03253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6023" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[8];
  assign _03255_ = _03254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6024" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[9];
  assign _03256_ = _03255_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6024" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[10];
  assign _03257_ = _03256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6025" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[11];
  assign _03258_ = _03257_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6025" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[12];
  assign _03259_ = _03258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6026" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[13];
  assign _03260_ = _03259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6026" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[14];
  assign _03261_ = _03260_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6027" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[15];
  assign _03262_ = _03261_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6027" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[16];
  assign _03263_ = _03262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6028" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[17];
  assign _03264_ = _03263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6028" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[18];
  assign _03265_ = _03264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6029" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[19];
  assign _03266_ = _03265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6029" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[20];
  assign _03267_ = _03266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6030" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[21];
  assign _03268_ = _03267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6030" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[22];
  assign _03269_ = _03268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6031" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[23];
  assign _03270_ = _03269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6031" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[24];
  assign _03271_ = _03270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6032" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[25];
  assign _03272_ = _03271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6032" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[26];
  assign _03273_ = _03272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6033" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[27];
  assign _03274_ = _03273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6033" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[28];
  assign _03275_ = _03274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6034" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[29];
  assign _03276_ = _03275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6034" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[30];
  assign _03277_ = _03276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6035" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[31];
  assign _03278_ = _03277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6035" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[32];
  assign _03279_ = _03278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6036" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[33];
  assign _03280_ = _03279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6036" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[34];
  assign _03281_ = _03280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6037" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[35];
  assign _03282_ = _03281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6037" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[36];
  assign _03283_ = _03282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6038" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[37];
  assign _03284_ = _03283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6038" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[38];
  assign _03285_ = _03284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6039" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[39];
  assign _03286_ = _03285_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6039" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[40];
  assign _03287_ = _03286_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6040" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[41];
  assign _03288_ = _03287_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6040" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[42];
  assign _03289_ = _03288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6041" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[43];
  assign _03290_ = _03289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6041" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[44];
  assign _03291_ = _03290_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6042" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[45];
  assign _03292_ = _03291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6042" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[46];
  assign _03293_ = _03292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6043" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[47];
  assign _03294_ = _03293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6043" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[48];
  assign _03295_ = _03294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6044" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[49];
  assign _03296_ = _03295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6044" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[50];
  assign _03297_ = _03296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6045" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[51];
  assign _03298_ = _03297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6045" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[52];
  assign _03299_ = _03298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6046" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[53];
  assign _03300_ = _03299_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6046" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[54];
  assign _03301_ = _03300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6047" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[55];
  assign _03302_ = _03301_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6047" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[56];
  assign _03303_ = _03302_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6048" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[57];
  assign _03304_ = _03303_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6048" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[58];
  assign _03305_ = _03304_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6049" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[59];
  assign _03306_ = _03305_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6049" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[60];
  assign _03307_ = _03306_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6050" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[61];
  assign _03308_ = _03307_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6050" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[62];
  assign _03309_ = _03308_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6051" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[63];
  assign _03310_ = _03309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6051" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[64];
  assign _03311_ = _03310_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6052" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[65];
  assign _03312_ = _03311_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6052" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[66];
  assign _03313_ = _03312_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6053" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[67];
  assign _03314_ = _03313_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6053" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[68];
  assign _03315_ = _03314_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6054" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[69];
  assign _03316_ = _03315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6054" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[70];
  assign _03317_ = _03316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6055" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[71];
  assign _03318_ = _03317_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6055" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[72];
  assign _03319_ = _03318_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6056" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[73];
  assign _03320_ = _03319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6056" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[74];
  assign _03321_ = _03320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6057" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[75];
  assign _03322_ = _03321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6057" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[76];
  assign _03323_ = _03322_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6058" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[77];
  assign _03324_ = _03323_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6058" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[78];
  assign _03325_ = _03324_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6059" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[79];
  assign _03326_ = _03325_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6059" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[80];
  assign _03327_ = _03326_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6060" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[81];
  assign _03328_ = _03327_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6060" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[82];
  assign _03329_ = _03328_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6061" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[83];
  assign _03330_ = _03329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6061" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[84];
  assign _03331_ = _03330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6062" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[85];
  assign _03332_ = _03331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6062" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[86];
  assign _03333_ = _03332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6063" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[87];
  assign _03334_ = _03333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6063" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[88];
  assign _03335_ = _03334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6064" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[89];
  assign _03336_ = _03335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6064" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[90];
  assign _03337_ = _03336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6065" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[91];
  assign _03338_ = _03337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6065" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[92];
  assign _03339_ = _03338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6066" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[93];
  assign _03340_ = _03339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6066" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[94];
  assign _03341_ = _03340_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6067" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[95];
  assign _03342_ = _03341_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6067" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[96];
  assign _03343_ = _03342_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6068" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[97];
  assign _03344_ = _03343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6068" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[98];
  assign _03345_ = _03344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6069" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[99];
  assign _03346_ = _03345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6069" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[100];
  assign _03347_ = _03346_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6070" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[101];
  assign _03348_ = _03347_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6070" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[102];
  assign _03349_ = _03348_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6071" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[103];
  assign _03350_ = _03349_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6071" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[104];
  assign _03351_ = _03350_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6072" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[105];
  assign _03352_ = _03351_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6072" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[106];
  assign _03353_ = _03352_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6073" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[107];
  assign _03354_ = _03353_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6073" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[108];
  assign _03355_ = _03354_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6074" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[109];
  assign _03356_ = _03355_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6074" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[110];
  assign _03357_ = _03356_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6075" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[111];
  assign _03358_ = _03357_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6075" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[112];
  assign _03359_ = _03358_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6076" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[113];
  assign _03360_ = _03359_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6076" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[114];
  assign _03361_ = _03360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6077" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[115];
  assign _03362_ = _03361_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6077" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[116];
  assign _03363_ = _03362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6078" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[117];
  assign _03364_ = _03363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6078" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[118];
  assign _03365_ = _03364_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6079" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[119];
  assign _03366_ = _03365_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6079" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[120];
  assign _03367_ = _03366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6080" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[121];
  assign _03368_ = _03367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6080" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[122];
  assign _03369_ = _03368_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6081" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[123];
  assign _03370_ = _03369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6081" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[124];
  assign _03371_ = _03370_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6082" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[125];
  assign _03372_ = _03371_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6082" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[126];
  assign _03373_ = _03372_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6083" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[127];
  assign _03374_ = _03373_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6083" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[128];
  assign _03375_ = _03374_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6084" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[129];
  assign _03376_ = _03375_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6084" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[130];
  assign _03377_ = _03376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6085" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[131];
  assign _03378_ = _03377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6085" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[132];
  assign _03379_ = _03378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6086" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[133];
  assign _03380_ = _03379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6086" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[134];
  assign _03381_ = _03380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6087" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[135];
  assign _03382_ = _03381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6087" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[136];
  assign _03383_ = _03382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6088" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[137];
  assign _03384_ = _03383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6088" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[138];
  assign _03385_ = _03384_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6089" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[139];
  assign _03386_ = _03385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6089" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[140];
  assign _03387_ = _03386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6090" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[141];
  assign _03388_ = _03387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6090" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[142];
  assign _03389_ = _03388_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6091" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[143];
  assign _03390_ = _03389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6091" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[144];
  assign _03391_ = _03390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6092" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[145];
  assign _03392_ = _03391_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6092" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[146];
  assign _03393_ = _03392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6093" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[147];
  assign _03394_ = _03393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6093" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[148];
  assign _03395_ = _03394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6094" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[149];
  assign _03396_ = _03395_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6094" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[150];
  assign _03397_ = _03396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6095" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[151];
  assign _03398_ = _03397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6095" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[152];
  assign _03399_ = _03398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6096" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[153];
  assign _03400_ = _03399_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6096" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[154];
  assign _03401_ = _03400_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6097" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[155];
  assign _03402_ = _03401_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6097" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[156];
  assign _03403_ = _03402_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6098" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[157];
  assign _03404_ = _03403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6098" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[158];
  assign _03405_ = _03404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6099" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[159];
  assign _03406_ = _03405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6099" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[160];
  assign _03407_ = _03406_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6100" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[161];
  assign _03408_ = _03407_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6100" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[162];
  assign _03409_ = _03408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6101" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[163];
  assign _03410_ = _03409_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6101" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[164];
  assign _03411_ = _03410_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6102" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[165];
  assign _03412_ = _03411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6102" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[166];
  assign _03413_ = _03412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6103" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[167];
  assign _03414_ = _03413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6103" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[168];
  assign _03415_ = _03414_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6104" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[169];
  assign _03416_ = _03415_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6104" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[170];
  assign _03417_ = _03416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6105" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[171];
  assign _03418_ = _03417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6105" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[172];
  assign _03419_ = _03418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6106" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[173];
  assign _03420_ = _03419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6106" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[174];
  assign _03421_ = _03420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6107" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[175];
  assign _03422_ = _03421_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6107" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[176];
  assign _03423_ = _03422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6108" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[177];
  assign _03424_ = _03423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6108" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[178];
  assign _03425_ = _03424_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6109" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[179];
  assign _03426_ = _03425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6109" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[180];
  assign _03427_ = _03426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6110" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[181];
  assign _03428_ = _03427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6110" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[182];
  assign _03429_ = _03428_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6111" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[183];
  assign _03430_ = _03429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6111" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[184];
  assign _03431_ = _03430_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6112" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[185];
  assign _03432_ = _03431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6112" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[186];
  assign _03433_ = _03432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6113" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[187];
  assign _03434_ = _03433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6113" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[188];
  assign _03435_ = _03434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6114" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[189];
  assign _03436_ = _03435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6114" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[190];
  assign _03437_ = _03436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6115" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[191];
  assign _03438_ = _03437_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6115" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[192];
  assign _03439_ = _03438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6116" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[193];
  assign _03440_ = _03439_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6116" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[194];
  assign _03441_ = _03440_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6117" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[195];
  assign _03442_ = _03441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6117" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[196];
  assign _03443_ = _03442_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6118" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[197];
  assign _03444_ = _03443_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6118" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[198];
  assign _03445_ = _03444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6119" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[199];
  assign _03446_ = _03445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6119" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[200];
  assign _03447_ = _03446_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6120" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[201];
  assign _03448_ = _03447_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6120" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[202];
  assign _03449_ = _03448_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6121" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[203];
  assign _03450_ = _03449_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6121" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[204];
  assign _03451_ = _03450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6122" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[205];
  assign _03452_ = _03451_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6122" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[206];
  assign _03453_ = _03452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6123" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[207];
  assign _03454_ = _03453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6123" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[208];
  assign _03455_ = _03454_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6124" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[209];
  assign _03456_ = _03455_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6124" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[210];
  assign _03457_ = _03456_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6125" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[211];
  assign _03458_ = _03457_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6125" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[212];
  assign _03459_ = _03458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6126" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[213];
  assign _03460_ = _03459_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6126" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[214];
  assign _03461_ = _03460_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6127" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[215];
  assign _03462_ = _03461_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6127" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[216];
  assign _03463_ = _03462_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6128" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[217];
  assign _03464_ = _03463_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6128" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[218];
  assign _03465_ = _03464_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6129" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[219];
  assign _03466_ = _03465_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6129" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[220];
  assign _03467_ = _03466_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6130" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[221];
  assign _03468_ = _03467_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6130" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[222];
  assign _03469_ = _03468_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6131" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[223];
  assign _03470_ = _03469_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6131" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[224];
  assign _03471_ = _03470_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6132" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[225];
  assign _03472_ = _03471_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6132" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[226];
  assign _03473_ = _03472_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6133" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[227];
  assign _03474_ = _03473_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6133" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[228];
  assign _03475_ = _03474_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6134" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[229];
  assign _03476_ = _03475_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6134" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[230];
  assign _03477_ = _03476_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6135" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[231];
  assign _03478_ = _03477_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6135" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[232];
  assign _03479_ = _03478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6136" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[233];
  assign _03480_ = _03479_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6136" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[234];
  assign _03481_ = _03480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6137" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[235];
  assign _03482_ = _03481_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6137" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[236];
  assign _03483_ = _03482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6138" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[237];
  assign _03484_ = _03483_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6138" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[238];
  assign _03485_ = _03484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6139" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[239];
  assign _03486_ = _03485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6139" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[240];
  assign _03487_ = _03486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6140" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[241];
  assign _03488_ = _03487_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6140" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[242];
  assign _03489_ = _03488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6141" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[243];
  assign _03490_ = _03489_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6141" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[244];
  assign _03491_ = _03490_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6142" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[245];
  assign _03492_ = _03491_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6142" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[246];
  assign _03493_ = _03492_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6143" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[247];
  assign _03494_ = _03493_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6143" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[248];
  assign _03495_ = _03494_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6144" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[249];
  assign _03496_ = _03495_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6144" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[250];
  assign _03497_ = _03496_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6145" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[251];
  assign _03498_ = _03497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6145" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[252];
  assign _03499_ = _03498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6146" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[253];
  assign _03500_ = _03499_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6146" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[254];
  assign _03501_ = _03500_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6147" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[255];
  assign _03502_ = _03501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6147" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[256];
  assign _03503_ = _03502_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6148" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[257];
  assign _03504_ = _03503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6148" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[258];
  assign _03505_ = _03504_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6149" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[259];
  assign _03506_ = _03505_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6149" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[260];
  assign _03507_ = _03506_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6150" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[261];
  assign _03508_ = _03507_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6150" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[262];
  assign _03509_ = _03508_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6151" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[263];
  assign _03510_ = _03509_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6151" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[264];
  assign _03511_ = _03510_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6152" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[265];
  assign _03512_ = _03511_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6152" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[266];
  assign _03513_ = _03512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6153" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[267];
  assign _03514_ = _03513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6153" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[268];
  assign _03515_ = _03514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6154" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[269];
  assign _03516_ = _03515_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6154" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[270];
  assign _03517_ = _03516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6155" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[271];
  assign _03518_ = _03517_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6155" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[272];
  assign _03519_ = _03518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6156" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[273];
  assign _03520_ = _03519_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6156" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[274];
  assign _03521_ = _03520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6157" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[275];
  assign _03522_ = _03521_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6157" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[276];
  assign _03523_ = _03522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6158" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[277];
  assign _03524_ = _03523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6158" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[278];
  assign _03525_ = _03524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6159" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[279];
  assign _03526_ = _03525_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6159" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[280];
  assign _03527_ = _03526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6160" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[281];
  assign _03528_ = _03527_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6160" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[282];
  assign _03529_ = _03528_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6161" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[283];
  assign _03530_ = _03529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6161" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[284];
  assign _03531_ = _03530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6162" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[285];
  assign _03532_ = _03531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6162" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[286];
  assign _03533_ = _03532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6163" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[287];
  assign _03534_ = _03533_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6163" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[288];
  assign _03535_ = _03534_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6164" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[289];
  assign _03536_ = _03535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6164" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[290];
  assign _03537_ = _03536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6165" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[291];
  assign _03538_ = _03537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6165" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[292];
  assign _03539_ = _03538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6166" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[293];
  assign _03540_ = _03539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6166" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[294];
  assign _03541_ = _03540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6167" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[295];
  assign _03542_ = _03541_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6167" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[296];
  assign _03543_ = _03542_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6168" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[297];
  assign _03544_ = _03543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6168" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[298];
  assign _03545_ = _03544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6169" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[299];
  assign _03546_ = _03545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6169" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[300];
  assign _03547_ = _03546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6170" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[301];
  assign _03548_ = _03547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6170" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[302];
  assign _03549_ = _03548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6171" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[303];
  assign _03550_ = _03549_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6171" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[304];
  assign _03551_ = _03550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6172" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[305];
  assign _03552_ = _03551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6172" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[306];
  assign _03553_ = _03552_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6173" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[307];
  assign _03554_ = _03553_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6173" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[308];
  assign _03555_ = _03554_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6174" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[309];
  assign _03556_ = _03555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6174" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[310];
  assign _03557_ = _03556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6175" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[311];
  assign _03558_ = _03557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6175" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[312];
  assign _03559_ = _03558_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6176" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[313];
  assign _03560_ = _03559_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6176" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[314];
  assign _03561_ = _03560_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6177" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[315];
  assign _03562_ = _03561_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6177" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[316];
  assign _03563_ = _03562_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6178" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[317];
  assign _03564_ = _03563_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6178" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[318];
  assign _03565_ = _03564_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6179" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[319];
  assign _03566_ = _03565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6179" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[320];
  assign _03567_ = _03566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6180" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[321];
  assign _03568_ = _03567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6180" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[322];
  assign _03569_ = _03568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6181" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[323];
  assign _03570_ = _03569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6181" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[324];
  assign _03571_ = _03570_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6182" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[325];
  assign _03572_ = _03571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6182" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[326];
  assign _03573_ = _03572_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6183" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[327];
  assign _03574_ = _03573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6183" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[328];
  assign _03575_ = _03574_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6184" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[329];
  assign _03576_ = _03575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6184" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[330];
  assign _03577_ = _03576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6185" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[331];
  assign _03578_ = _03577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6185" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[332];
  assign _03579_ = _03578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6186" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[333];
  assign _03580_ = _03579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6186" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[334];
  assign _03581_ = _03580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6187" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[335];
  assign _03582_ = _03581_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6187" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[336];
  assign _03583_ = _03582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6188" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[337];
  assign _03584_ = _03583_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6188" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[338];
  assign _03585_ = _03584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6189" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[339];
  assign _03586_ = _03585_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6189" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[340];
  assign _03587_ = _03586_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6190" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[341];
  assign _03588_ = _03587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6190" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[342];
  assign _03589_ = _03588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6191" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[343];
  assign _03590_ = _03589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6191" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[344];
  assign _03591_ = _03590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6192" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[345];
  assign _03592_ = _03591_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6192" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[346];
  assign _03593_ = _03592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6193" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[347];
  assign _03594_ = _03593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6193" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[348];
  assign _03595_ = _03594_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6194" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[349];
  assign _03596_ = _03595_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6194" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[350];
  assign _03597_ = _03596_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6195" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[351];
  assign _03598_ = _03597_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6195" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[352];
  assign _03599_ = _03598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6196" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[353];
  assign _03600_ = _03599_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6196" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[354];
  assign _03601_ = _03600_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6197" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[355];
  assign _03602_ = _03601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6197" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[356];
  assign _03603_ = _03602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6198" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[357];
  assign _03604_ = _03603_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6198" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[358];
  assign _03605_ = _03604_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6199" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[359];
  assign _03606_ = _03605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6199" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[360];
  assign _03607_ = _03606_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6200" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[361];
  assign _03608_ = _03607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6200" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[362];
  assign _03609_ = _03608_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6201" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[363];
  assign _03610_ = _03609_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6201" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[364];
  assign _03611_ = _03610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6202" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[365];
  assign _03612_ = _03611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6202" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[366];
  assign _03613_ = _03612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6203" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[367];
  assign _03614_ = _03613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6203" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[368];
  assign _03615_ = _03614_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6204" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[369];
  assign _03616_ = _03615_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6204" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[370];
  assign _03617_ = _03616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6205" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[371];
  assign _03618_ = _03617_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6205" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[372];
  assign _03619_ = _03618_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6206" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[373];
  assign _03620_ = _03619_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6206" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[374];
  assign _03621_ = _03620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6207" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[375];
  assign _03622_ = _03621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6207" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[376];
  assign _03623_ = _03622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6208" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[377];
  assign _03624_ = _03623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6208" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[378];
  assign _03625_ = _03624_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6209" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[379];
  assign _03626_ = _03625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6209" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[380];
  assign _03627_ = _03626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6210" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[381];
  assign _03628_ = _03627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6210" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[382];
  assign _03629_ = _03628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6211" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[383];
  assign _03630_ = _03629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6211" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[384];
  assign _03631_ = _03630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6212" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[385];
  assign _03632_ = _03631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6212" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[386];
  assign _03633_ = _03632_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6213" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[387];
  assign _03634_ = _03633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6213" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[388];
  assign _03635_ = _03634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6214" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[389];
  assign _03636_ = _03635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6214" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[390];
  assign _03637_ = _03636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6215" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[391];
  assign _03638_ = _03637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6215" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[392];
  assign _03639_ = _03638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6216" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[393];
  assign _03640_ = _03639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6216" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[394];
  assign _03641_ = _03640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6217" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[395];
  assign _03642_ = _03641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6217" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[396];
  assign _03643_ = _03642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6218" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[397];
  assign _03644_ = _03643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6218" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[398];
  assign _03645_ = _03644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6219" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[399];
  assign _03646_ = _03645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6219" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[400];
  assign _03647_ = _03646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6220" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[401];
  assign _03648_ = _03647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6220" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[402];
  assign _03649_ = _03648_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6221" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[403];
  assign _03650_ = _03649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6221" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[404];
  assign _03651_ = _03650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6222" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[405];
  assign _03652_ = _03651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6222" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[406];
  assign _03653_ = _03652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6223" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[407];
  assign _03654_ = _03653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6223" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[408];
  assign _03655_ = _03654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6224" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[409];
  assign _03656_ = _03655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6224" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[410];
  assign _03657_ = _03656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6225" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[411];
  assign _03658_ = _03657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6225" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[412];
  assign _03659_ = _03658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6226" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[413];
  assign _03660_ = _03659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6226" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[414];
  assign _03661_ = _03660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6227" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[415];
  assign _03662_ = _03661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6227" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[416];
  assign _03663_ = _03662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6228" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[417];
  assign _03664_ = _03663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6228" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[418];
  assign _03665_ = _03664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6229" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[419];
  assign _03666_ = _03665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6229" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[420];
  assign _03667_ = _03666_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6230" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[421];
  assign _03668_ = _03667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6230" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[422];
  assign _03669_ = _03668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6231" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[423];
  assign _03670_ = _03669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6231" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[424];
  assign _03671_ = _03670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6232" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[425];
  assign _03672_ = _03671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6232" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[426];
  assign _03673_ = _03672_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6233" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[427];
  assign _03674_ = _03673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6233" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[428];
  assign _03675_ = _03674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6234" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[429];
  assign _03676_ = _03675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6234" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[430];
  assign _03677_ = _03676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6235" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[431];
  assign _03678_ = _03677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6235" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[432];
  assign _03679_ = _03678_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6236" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[433];
  assign _03680_ = _03679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6236" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[434];
  assign _03681_ = _03680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6237" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[435];
  assign _03682_ = _03681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6237" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[436];
  assign _03683_ = _03682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6238" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[437];
  assign _03684_ = _03683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6238" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[438];
  assign _03685_ = _03684_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6239" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[439];
  assign _03686_ = _03685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6239" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[440];
  assign _03687_ = _03686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6240" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[441];
  assign _03688_ = _03687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6240" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[442];
  assign _03689_ = _03688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6241" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[443];
  assign _03690_ = _03689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6241" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[444];
  assign _03691_ = _03690_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6242" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[445];
  assign _03692_ = _03691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6242" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[446];
  assign _03693_ = _03692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6243" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[447];
  assign _03694_ = _03693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6243" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[448];
  assign _03695_ = _03694_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6244" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[449];
  assign _03696_ = _03695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6244" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[450];
  assign _03697_ = _03696_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6245" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[451];
  assign _03698_ = _03697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6245" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[452];
  assign _03699_ = _03698_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6246" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[453];
  assign _03700_ = _03699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6246" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[454];
  assign _03701_ = _03700_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6247" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[455];
  assign _03702_ = _03701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6247" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[456];
  assign _03703_ = _03702_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6248" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[457];
  assign _03704_ = _03703_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6248" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[458];
  assign _03705_ = _03704_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6249" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[459];
  assign _03706_ = _03705_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6249" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[460];
  assign _03707_ = _03706_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6250" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[461];
  assign _03708_ = _03707_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6250" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[462];
  assign _03709_ = _03708_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6251" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[463];
  assign _03710_ = _03709_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6251" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[464];
  assign _03711_ = _03710_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6252" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[465];
  assign _03712_ = _03711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6252" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[466];
  assign _03713_ = _03712_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6253" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[467];
  assign _03714_ = _03713_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6253" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[468];
  assign _03715_ = _03714_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6254" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[469];
  assign _03716_ = _03715_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6254" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[470];
  assign _03717_ = _03716_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6255" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[471];
  assign _03718_ = _03717_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6255" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[472];
  assign _03719_ = _03718_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6256" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[473];
  assign _03720_ = _03719_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6256" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[474];
  assign _03721_ = _03720_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6257" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[475];
  assign _03722_ = _03721_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6257" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[476];
  assign _03723_ = _03722_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6258" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[477];
  assign _03724_ = _03723_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6258" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[478];
  assign _03725_ = _03724_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6259" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[479];
  assign _03726_ = _03725_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6259" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[480];
  assign _03727_ = _03726_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6260" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[481];
  assign _03728_ = _03727_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6260" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[482];
  assign _03729_ = _03728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6261" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[483];
  assign _03730_ = _03729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6261" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[484];
  assign _03731_ = _03730_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6262" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[485];
  assign _03732_ = _03731_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6262" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[486];
  assign _03733_ = _03732_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6263" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[487];
  assign _03734_ = _03733_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6263" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[488];
  assign _03735_ = _03734_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6264" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[489];
  assign _03736_ = _03735_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6264" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[490];
  assign _03737_ = _03736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6265" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[491];
  assign _03738_ = _03737_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6265" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[492];
  assign _03739_ = _03738_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6266" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[493];
  assign _03740_ = _03739_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6266" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[494];
  assign _03741_ = _03740_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6267" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[495];
  assign _03742_ = _03741_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6267" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[496];
  assign _03743_ = _03742_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6268" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[497];
  assign _03744_ = _03743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6268" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[498];
  assign _03745_ = _03744_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6269" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[499];
  assign _03746_ = _03745_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6269" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[500];
  assign _03747_ = _03746_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6270" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[501];
  assign _03748_ = _03747_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6270" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[502];
  assign _03749_ = _03748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6271" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[503];
  assign _03750_ = _03749_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6271" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[504];
  assign _03751_ = _03750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6272" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[505];
  assign _03752_ = _03751_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6272" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[506];
  assign _03753_ = _03752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6273" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[507];
  assign _03754_ = _03753_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6273" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[508];
  assign _03755_ = _03754_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6274" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[509];
  assign _03756_ = _03755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6274" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[510];
  assign _03757_ = _03756_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6275" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[511];
  assign _03758_ = _03757_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6275" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[512];
  assign _03759_ = _03758_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6276" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[513];
  assign _03760_ = _03759_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6276" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[514];
  assign _03761_ = _03760_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6277" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[515];
  assign _03762_ = _03761_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6277" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[516];
  assign _03763_ = _03762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6278" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[517];
  assign _03764_ = _03763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6278" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[518];
  assign _03765_ = _03764_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6279" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[519];
  assign _03766_ = _03765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6279" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[520];
  assign _03767_ = _03766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6280" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[521];
  assign _03768_ = _03767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6280" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[522];
  assign _03769_ = _03768_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6281" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[523];
  assign _03770_ = _03769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6281" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[524];
  assign _03771_ = _03770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6282" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[525];
  assign _03772_ = _03771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6282" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[526];
  assign _03773_ = _03772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6283" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[527];
  assign _03774_ = _03773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6283" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[528];
  assign _03775_ = _03774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6284" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[529];
  assign _03776_ = _03775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6284" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[530];
  assign _03777_ = _03776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6285" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[531];
  assign _03778_ = _03777_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6285" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[532];
  assign _03779_ = _03778_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6286" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[533];
  assign _03780_ = _03779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6286" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[534];
  assign _03781_ = _03780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6287" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[535];
  assign _03782_ = _03781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6287" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[536];
  assign _03783_ = _03782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6288" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[537];
  assign _03784_ = _03783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6288" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[538];
  assign _03785_ = _03784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6289" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[539];
  assign _03786_ = _03785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6289" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[540];
  assign _03787_ = _03786_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6290" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[541];
  assign _03788_ = _03787_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6290" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[542];
  assign _03789_ = _03788_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6291" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[543];
  assign _03790_ = _03789_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6291" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[544];
  assign _03791_ = _03790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6292" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[545];
  assign _03792_ = _03791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6292" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[546];
  assign _03793_ = _03792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6293" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[547];
  assign _03794_ = _03793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6293" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[548];
  assign _03795_ = _03794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6294" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[549];
  assign _03796_ = _03795_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6294" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[550];
  assign _03797_ = _03796_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6295" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[551];
  assign _03798_ = _03797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6295" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[552];
  assign _03799_ = _03798_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6296" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[553];
  assign _03800_ = _03799_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6296" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[554];
  assign _03801_ = _03800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6297" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[555];
  assign _03802_ = _03801_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6297" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[556];
  assign _03803_ = _03802_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6298" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[557];
  assign _03804_ = _03803_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6298" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[558];
  assign _03805_ = _03804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6299" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[559];
  assign _03806_ = _03805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6299" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[560];
  assign _03807_ = _03806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6300" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[561];
  assign _03808_ = _03807_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6300" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[562];
  assign _03809_ = _03808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6301" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[563];
  assign _03810_ = _03809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6301" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[564];
  assign _03811_ = _03810_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6302" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[565];
  assign _03812_ = _03811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6302" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[566];
  assign _03813_ = _03812_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6303" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[567];
  assign _03814_ = _03813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6303" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[568];
  assign _03815_ = _03814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6304" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[569];
  assign _03816_ = _03815_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6304" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[570];
  assign _03817_ = _03816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6305" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[571];
  assign _03818_ = _03817_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6305" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[572];
  assign _03819_ = _03818_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6306" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[573];
  assign _03820_ = _03819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6306" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[574];
  assign _03821_ = _03820_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6307" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[575];
  assign _03822_ = _03821_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6307" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[576];
  assign _03823_ = _03822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6308" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[577];
  assign _03824_ = _03823_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6308" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[578];
  assign _03825_ = _03824_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6309" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[579];
  assign _03826_ = _03825_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6309" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[580];
  assign _03827_ = _03826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6310" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[581];
  assign _03828_ = _03827_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6310" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[582];
  assign _03829_ = _03828_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6311" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[583];
  assign _03830_ = _03829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6311" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[584];
  assign _03831_ = _03830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6312" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[585];
  assign _03832_ = _03831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6312" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[586];
  assign _03833_ = _03832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6313" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[587];
  assign _03834_ = _03833_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6313" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[588];
  assign _03835_ = _03834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6314" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[589];
  assign _03836_ = _03835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6314" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[590];
  assign _03837_ = _03836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6315" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[591];
  assign _03838_ = _03837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6315" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[592];
  assign _03839_ = _03838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6316" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[593];
  assign _03840_ = _03839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6316" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[594];
  assign _03841_ = _03840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6317" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[595];
  assign _03842_ = _03841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6317" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[596];
  assign _03843_ = _03842_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6318" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[597];
  assign _03844_ = _03843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6318" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[598];
  assign _03845_ = _03844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6319" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[599];
  assign _03846_ = _03845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6319" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[600];
  assign _03847_ = _03846_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6320" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[601];
  assign _03848_ = _03847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6320" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[602];
  assign _03849_ = _03848_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6321" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[603];
  assign _03850_ = _03849_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6321" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[604];
  assign _03851_ = _03850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6322" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[605];
  assign _03852_ = _03851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6322" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[606];
  assign _03853_ = _03852_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6323" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[607];
  assign _03854_ = _03853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6323" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[608];
  assign _03855_ = _03854_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6324" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[609];
  assign _03856_ = _03855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6324" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[610];
  assign _03857_ = _03856_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6325" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[611];
  assign _03858_ = _03857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6325" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[612];
  assign _03859_ = _03858_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6326" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[613];
  assign _03860_ = _03859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6326" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[614];
  assign _03861_ = _03860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6327" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[615];
  assign _03862_ = _03861_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6327" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[616];
  assign _03863_ = _03862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6328" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[617];
  assign _03864_ = _03863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6328" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[618];
  assign _03865_ = _03864_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6329" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[619];
  assign _03866_ = _03865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6329" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[620];
  assign _03867_ = _03866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6330" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[621];
  assign _03868_ = _03867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6330" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[622];
  assign _03869_ = _03868_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6331" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[623];
  assign _03870_ = _03869_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6331" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[624];
  assign _03871_ = _03870_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6332" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[625];
  assign _03872_ = _03871_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6332" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[626];
  assign _03873_ = _03872_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6333" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[627];
  assign _03874_ = _03873_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6333" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[628];
  assign _03875_ = _03874_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6334" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[629];
  assign _03876_ = _03875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6334" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[630];
  assign _03877_ = _03876_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6335" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[631];
  assign _03878_ = _03877_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6335" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[632];
  assign _03879_ = _03878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6336" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[633];
  assign _03880_ = _03879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6336" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[634];
  assign _03881_ = _03880_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6337" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[635];
  assign _03882_ = _03881_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6337" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[636];
  assign _03883_ = _03882_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6338" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[637];
  assign _03884_ = _03883_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6338" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[638];
  assign _03885_ = _03884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6339" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[639];
  assign _03886_ = _03885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6339" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[640];
  assign _03887_ = _03886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6340" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[641];
  assign _03888_ = _03887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6340" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[642];
  assign _03889_ = _03888_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6341" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[643];
  assign _03890_ = _03889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6341" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[644];
  assign _03891_ = _03890_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6342" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[645];
  assign _03892_ = _03891_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6342" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[646];
  assign _03893_ = _03892_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6343" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[647];
  assign _03894_ = _03893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6343" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[648];
  assign _03895_ = _03894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6344" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[649];
  assign _03896_ = _03895_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6344" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[650];
  assign _03897_ = _03896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6345" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[651];
  assign _03898_ = _03897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6345" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[652];
  assign _03899_ = _03898_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6346" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[653];
  assign _03900_ = _03899_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6346" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[654];
  assign _03901_ = _03900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6347" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[655];
  assign _03902_ = _03901_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6347" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[656];
  assign _03903_ = _03902_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6348" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[657];
  assign _03904_ = _03903_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6348" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[658];
  assign _03905_ = _03904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6349" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[659];
  assign _03906_ = _03905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6349" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[660];
  assign _03907_ = _03906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6350" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[661];
  assign _03908_ = _03907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6350" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[662];
  assign _03909_ = _03908_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6351" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[663];
  assign _03910_ = _03909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6351" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[664];
  assign _03911_ = _03910_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6352" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[665];
  assign _03912_ = _03911_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6352" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[666];
  assign _03913_ = _03912_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6353" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[667];
  assign _03914_ = _03913_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6353" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[668];
  assign _03915_ = _03914_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6354" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[669];
  assign _03916_ = _03915_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6354" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[670];
  assign _03917_ = _03916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6355" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[671];
  assign _03918_ = _03917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6355" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[672];
  assign _03919_ = _03918_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6356" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[673];
  assign _03920_ = _03919_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6356" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[674];
  assign _03921_ = _03920_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6357" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[675];
  assign _03922_ = _03921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6357" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[676];
  assign _03923_ = _03922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6358" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[677];
  assign _03924_ = _03923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6358" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[678];
  assign _03925_ = _03924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6359" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[679];
  assign _03926_ = _03925_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6359" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[680];
  assign _03927_ = _03926_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6360" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[681];
  assign _03928_ = _03927_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6360" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[682];
  assign _03929_ = _03928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6361" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[683];
  assign _03930_ = _03929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6361" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[684];
  assign _03931_ = _03930_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6362" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[685];
  assign _03932_ = _03931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6362" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[686];
  assign _03933_ = _03932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6363" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[687];
  assign _03934_ = _03933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6363" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[688];
  assign _03935_ = _03934_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6364" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[689];
  assign _03936_ = _03935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6364" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[690];
  assign _03937_ = _03936_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6365" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[691];
  assign _03938_ = _03937_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6365" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[692];
  assign _03939_ = _03938_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6366" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[693];
  assign _03940_ = _03939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6366" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[694];
  assign _03941_ = _03940_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6367" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[695];
  assign _03942_ = _03941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6367" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[696];
  assign _03943_ = _03942_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6368" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[697];
  assign _03944_ = _03943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6368" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[698];
  assign _03945_ = _03944_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6369" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[699];
  assign _03946_ = _03945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6369" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[700];
  assign _03947_ = _03946_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6370" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[701];
  assign _03948_ = _03947_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6370" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[702];
  assign _03949_ = _03948_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6371" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[703];
  assign _03950_ = _03949_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6371" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[704];
  assign _03951_ = _03950_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6372" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[705];
  assign _03952_ = _03951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6372" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[706];
  assign _03953_ = _03952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6373" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[707];
  assign _03954_ = _03953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6373" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[708];
  assign _03955_ = _03954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6374" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[709];
  assign _03956_ = _03955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6374" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[710];
  assign _03957_ = _03956_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6375" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[711];
  assign _03958_ = _03957_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6375" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[712];
  assign _03959_ = _03958_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6376" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[713];
  assign _03960_ = _03959_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6376" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[714];
  assign _03961_ = _03960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6377" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[715];
  assign _03962_ = _03961_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6377" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[716];
  assign _03963_ = _03962_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6378" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[717];
  assign _03964_ = _03963_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6378" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[718];
  assign _03965_ = _03964_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6379" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[719];
  assign _03966_ = _03965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6379" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[720];
  assign _03967_ = _03966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6380" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[721];
  assign _03968_ = _03967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6380" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[722];
  assign _03969_ = _03968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6381" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[723];
  assign _03970_ = _03969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6381" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[724];
  assign _03971_ = _03970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6382" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[725];
  assign _03972_ = _03971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6382" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[726];
  assign _03973_ = _03972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6383" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[727];
  assign _03974_ = _03973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6383" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[728];
  assign _03975_ = _03974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6384" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[729];
  assign _03976_ = _03975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6384" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[730];
  assign _03977_ = _03976_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6385" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[731];
  assign _03978_ = _03977_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6385" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[732];
  assign _03979_ = _03978_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6386" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[733];
  assign _03980_ = _03979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6386" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[734];
  assign _03981_ = _03980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6387" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[735];
  assign _03982_ = _03981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6387" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[736];
  assign _03983_ = _03982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6388" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[737];
  assign _03984_ = _03983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6388" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[738];
  assign _03985_ = _03984_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6389" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[739];
  assign _03986_ = _03985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6389" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[740];
  assign _03987_ = _03986_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6390" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[741];
  assign _03988_ = _03987_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6390" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[742];
  assign _03989_ = _03988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6391" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[743];
  assign _03990_ = _03989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6391" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[744];
  assign _03991_ = _03990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6392" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[745];
  assign _03992_ = _03991_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6392" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[746];
  assign _03993_ = _03992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6393" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[747];
  assign _03994_ = _03993_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6393" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[748];
  assign _03995_ = _03994_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6394" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[749];
  assign _03996_ = _03995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6394" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[750];
  assign _03997_ = _03996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6395" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[751];
  assign _03998_ = _03997_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6395" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[752];
  assign _03999_ = _03998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6396" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[753];
  assign _04000_ = _03999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6396" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[754];
  assign _04001_ = _04000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6397" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[755];
  assign _04002_ = _04001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6397" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[756];
  assign _04003_ = _04002_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6398" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[757];
  assign _04004_ = _04003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6398" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[758];
  assign _04005_ = _04004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6399" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[759];
  assign _04006_ = _04005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6399" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[760];
  assign _04007_ = _04006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6400" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[761];
  assign _04008_ = _04007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6400" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[762];
  assign _04009_ = _04008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6401" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[763];
  assign _04010_ = _04009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6401" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[764];
  assign _04011_ = _04010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6402" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[765];
  assign _04012_ = _04011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6402" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[766];
  assign _04013_ = _04012_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6403" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[767];
  assign _04014_ = _04013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6403" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[768];
  assign _04015_ = _04014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6404" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[769];
  assign _04016_ = _04015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6404" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[770];
  assign _04017_ = _04016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6405" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[771];
  assign _04018_ = _04017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6405" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[772];
  assign _04019_ = _04018_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6406" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[773];
  assign _04020_ = _04019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6406" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[774];
  assign _04021_ = _04020_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6407" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[775];
  assign _04022_ = _04021_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6407" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[776];
  assign _04023_ = _04022_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6408" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[777];
  assign _04024_ = _04023_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6408" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[778];
  assign _04025_ = _04024_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6409" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[779];
  assign _04026_ = _04025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6409" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[780];
  assign _04027_ = _04026_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6410" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[781];
  assign _04028_ = _04027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6410" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[782];
  assign _04029_ = _04028_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6411" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[783];
  assign _04030_ = _04029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6411" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[784];
  assign _04031_ = _04030_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6412" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[785];
  assign _04032_ = _04031_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6412" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[786];
  assign _04033_ = _04032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6413" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[787];
  assign _04034_ = _04033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6413" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[788];
  assign _04035_ = _04034_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6414" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[789];
  assign _04036_ = _04035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6414" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[790];
  assign _04037_ = _04036_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6415" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[791];
  assign _04038_ = _04037_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6415" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[792];
  assign _04039_ = _04038_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6416" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[793];
  assign _04040_ = _04039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6416" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[794];
  assign _04041_ = _04040_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6417" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[795];
  assign _04042_ = _04041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6417" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[796];
  assign _04043_ = _04042_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6418" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[797];
  assign _04044_ = _04043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6418" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[798];
  assign _04045_ = _04044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6419" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[799];
  assign _04046_ = _04045_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6419" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[800];
  assign _04047_ = _04046_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6420" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[801];
  assign _04048_ = _04047_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6420" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[802];
  assign _04049_ = _04048_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6421" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[803];
  assign _04050_ = _04049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6421" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[804];
  assign _04051_ = _04050_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6422" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[805];
  assign _04052_ = _04051_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6422" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[806];
  assign _04053_ = _04052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6423" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[807];
  assign _04054_ = _04053_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6423" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[808];
  assign _04055_ = _04054_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6424" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[809];
  assign _04056_ = _04055_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6424" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[810];
  assign _04057_ = _04056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6425" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[811];
  assign _04058_ = _04057_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6425" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[812];
  assign _04059_ = _04058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6426" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[813];
  assign _04060_ = _04059_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6426" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[814];
  assign _04061_ = _04060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6427" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[815];
  assign _04062_ = _04061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6427" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[816];
  assign _04063_ = _04062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6428" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[817];
  assign _04064_ = _04063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6428" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[818];
  assign _04065_ = _04064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6429" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[819];
  assign _04066_ = _04065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6429" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[820];
  assign _04067_ = _04066_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6430" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[821];
  assign _04068_ = _04067_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6430" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[822];
  assign _04069_ = _04068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6431" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[823];
  assign _04070_ = _04069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6431" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[824];
  assign _04071_ = _04070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6432" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[825];
  assign _04072_ = _04071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6432" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[826];
  assign _04073_ = _04072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6433" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[827];
  assign _04074_ = _04073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6433" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[828];
  assign _04075_ = _04074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6434" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[829];
  assign _04076_ = _04075_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6434" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[830];
  assign _04077_ = _04076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6435" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[831];
  assign _04078_ = _04077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6435" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[832];
  assign _04079_ = _04078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6436" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[833];
  assign _04080_ = _04079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6436" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[834];
  assign _04081_ = _04080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6437" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[835];
  assign _04082_ = _04081_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6437" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[836];
  assign _04083_ = _04082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6438" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[837];
  assign _04084_ = _04083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6438" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[838];
  assign _04085_ = _04084_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6439" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[839];
  assign _04086_ = _04085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6439" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[840];
  assign _04087_ = _04086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6440" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[841];
  assign _04088_ = _04087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6440" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[842];
  assign _04089_ = _04088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6441" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[843];
  assign _04090_ = _04089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6441" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[844];
  assign _04091_ = _04090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6442" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[845];
  assign _04092_ = _04091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6442" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[846];
  assign _04093_ = _04092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6443" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[847];
  assign _04094_ = _04093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6443" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[848];
  assign _04095_ = _04094_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6444" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[849];
  assign _04096_ = _04095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6444" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[850];
  assign _04097_ = _04096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6445" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[851];
  assign _04098_ = _04097_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6445" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[852];
  assign _04099_ = _04098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6446" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[853];
  assign _04100_ = _04099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6446" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[854];
  assign _04101_ = _04100_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6447" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[855];
  assign _04102_ = _04101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6447" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[856];
  assign _04103_ = _04102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6448" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[857];
  assign _04104_ = _04103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6448" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[858];
  assign _04105_ = _04104_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6449" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[859];
  assign _04106_ = _04105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6449" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[860];
  assign _04107_ = _04106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6450" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[861];
  assign _04108_ = _04107_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6450" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[862];
  assign _04109_ = _04108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6451" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[863];
  assign _04110_ = _04109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6451" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[864];
  assign _04111_ = _04110_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6452" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[865];
  assign _04112_ = _04111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6452" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[866];
  assign _04113_ = _04112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6453" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[867];
  assign _04114_ = _04113_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6453" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[868];
  assign _04115_ = _04114_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6454" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[869];
  assign _04116_ = _04115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6454" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[870];
  assign _04117_ = _04116_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6455" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[871];
  assign _04118_ = _04117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6455" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[872];
  assign _04119_ = _04118_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6456" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[873];
  assign _04120_ = _04119_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6456" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[874];
  assign _04121_ = _04120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6457" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[875];
  assign _04122_ = _04121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6457" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[876];
  assign _04123_ = _04122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6458" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[877];
  assign _04124_ = _04123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6458" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[878];
  assign _04125_ = _04124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6459" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[879];
  assign _04126_ = _04125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6459" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[880];
  assign _04127_ = _04126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6460" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[881];
  assign _04128_ = _04127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6460" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[882];
  assign _04129_ = _04128_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6461" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[883];
  assign _04130_ = _04129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6461" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[884];
  assign _04131_ = _04130_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6462" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[885];
  assign _04132_ = _04131_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6462" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[886];
  assign _04133_ = _04132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6463" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[887];
  assign _04134_ = _04133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6463" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[888];
  assign _04135_ = _04134_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6464" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[889];
  assign _04136_ = _04135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6464" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[890];
  assign _04137_ = _04136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6465" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[891];
  assign _04138_ = _04137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6465" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[892];
  assign _04139_ = _04138_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6466" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[893];
  assign _04140_ = _04139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6466" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[894];
  assign _04141_ = _04140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6467" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[895];
  assign _04142_ = _04141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6467" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[896];
  assign _04143_ = _04142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6468" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[897];
  assign _04144_ = _04143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6468" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[898];
  assign _04145_ = _04144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6469" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[899];
  assign _04146_ = _04145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6469" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[900];
  assign _04147_ = _04146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6470" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[901];
  assign _04148_ = _04147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6470" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[902];
  assign _04149_ = _04148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6471" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[903];
  assign _04150_ = _04149_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6471" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[904];
  assign _04151_ = _04150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6472" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[905];
  assign _04152_ = _04151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6472" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[906];
  assign _04153_ = _04152_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6473" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[907];
  assign _04154_ = _04153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6473" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[908];
  assign _04155_ = _04154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6474" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[909];
  assign _04156_ = _04155_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6474" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[910];
  assign _04157_ = _04156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6475" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[911];
  assign _04158_ = _04157_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6475" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[912];
  assign _04159_ = _04158_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6476" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[913];
  assign _04160_ = _04159_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6476" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[914];
  assign _04161_ = _04160_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6477" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[915];
  assign _04162_ = _04161_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6477" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[916];
  assign _04163_ = _04162_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6478" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[917];
  assign _04164_ = _04163_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6478" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[918];
  assign _04165_ = _04164_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6479" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[919];
  assign _04166_ = _04165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6479" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[920];
  assign _04167_ = _04166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6480" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[921];
  assign _04168_ = _04167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6480" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[922];
  assign _04169_ = _04168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6481" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[923];
  assign _04170_ = _04169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6481" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[924];
  assign _04171_ = _04170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6482" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[925];
  assign _04172_ = _04171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6482" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[926];
  assign _04173_ = _04172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6483" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[927];
  assign _04174_ = _04173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6483" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[928];
  assign _04175_ = _04174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6484" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[929];
  assign _04176_ = _04175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6484" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[930];
  assign _04177_ = _04176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6485" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[931];
  assign _04178_ = _04177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6485" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[932];
  assign _04179_ = _04178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6486" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[933];
  assign _04180_ = _04179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6486" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[934];
  assign _04181_ = _04180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6487" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[935];
  assign _04182_ = _04181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6487" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[936];
  assign _04183_ = _04182_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6488" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[937];
  assign _04184_ = _04183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6488" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[938];
  assign _04185_ = _04184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6489" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[939];
  assign _04186_ = _04185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6489" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[940];
  assign _04187_ = _04186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6490" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[941];
  assign _04188_ = _04187_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6490" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[942];
  assign _04189_ = _04188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6491" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[943];
  assign _04190_ = _04189_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6491" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[944];
  assign _04191_ = _04190_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6492" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[945];
  assign _04192_ = _04191_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6492" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[946];
  assign _04193_ = _04192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6493" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[947];
  assign _04194_ = _04193_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6493" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[948];
  assign _04195_ = _04194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6494" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[949];
  assign _04196_ = _04195_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6494" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[950];
  assign _04197_ = _04196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6495" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[951];
  assign _04198_ = _04197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6495" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[952];
  assign _04199_ = _04198_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6496" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[953];
  assign _04200_ = _04199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6496" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[954];
  assign _04201_ = _04200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6497" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[955];
  assign _04202_ = _04201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6497" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[956];
  assign _04203_ = _04202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6498" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[957];
  assign _04204_ = _04203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6498" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[958];
  assign _04205_ = _04204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6499" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[959];
  assign _04206_ = _04205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6499" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[960];
  assign _04207_ = _04206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6500" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[961];
  assign _04208_ = _04207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6500" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[962];
  assign _04209_ = _04208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6501" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[963];
  assign _04210_ = _04209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6501" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[964];
  assign _04211_ = _04210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6502" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[965];
  assign _04212_ = _04211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6502" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[966];
  assign _04213_ = _04212_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6503" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[967];
  assign _04214_ = _04213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6503" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[968];
  assign _04215_ = _04214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6504" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[969];
  assign _04216_ = _04215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6504" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[970];
  assign _04217_ = _04216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6505" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[971];
  assign _04218_ = _04217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6505" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[972];
  assign _04219_ = _04218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6506" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[973];
  assign _04220_ = _04219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6506" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[974];
  assign _04221_ = _04220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6507" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[975];
  assign _04222_ = _04221_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6507" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[976];
  assign _04223_ = _04222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6508" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[977];
  assign _04224_ = _04223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6508" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[978];
  assign _04225_ = _04224_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6509" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[979];
  assign _04226_ = _04225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6509" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[980];
  assign _04227_ = _04226_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6510" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[981];
  assign _04228_ = _04227_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6510" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[982];
  assign _04229_ = _04228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6511" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[983];
  assign _04230_ = _04229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6511" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[984];
  assign _04231_ = _04230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6512" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[985];
  assign _04232_ = _04231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6512" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[986];
  assign _04233_ = _04232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6513" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[987];
  assign _04234_ = _04233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6513" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[988];
  assign _04235_ = _04234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6514" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[989];
  assign _04236_ = _04235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6514" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[990];
  assign _04237_ = _04236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6515" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[991];
  assign _04238_ = _04237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6515" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[992];
  assign _04239_ = _04238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6516" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[993];
  assign _04240_ = _04239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6516" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[994];
  assign _04241_ = _04240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6517" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[995];
  assign _04242_ = _04241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6517" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[996];
  assign _04243_ = _04242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6518" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[997];
  assign _04244_ = _04243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6518" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[998];
  assign _04245_ = _04244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6519" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[999];
  assign _04246_ = _04245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6519" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1000];
  assign _04247_ = _04246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6520" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1001];
  assign _04248_ = _04247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6520" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1002];
  assign _04249_ = _04248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6521" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1003];
  assign _04250_ = _04249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6521" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1004];
  assign _04251_ = _04250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6522" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1005];
  assign _04252_ = _04251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6522" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1006];
  assign _04253_ = _04252_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6523" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1007];
  assign _04254_ = _04253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6523" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1008];
  assign _04255_ = _04254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6524" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1009];
  assign _04256_ = _04255_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6524" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1010];
  assign _04257_ = _04256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6525" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1011];
  assign _04258_ = _04257_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6525" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1012];
  assign _04259_ = _04258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6526" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1013];
  assign _04260_ = _04259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6526" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1014];
  assign _04261_ = _04260_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6527" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1015];
  assign _04262_ = _04261_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6527" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1016];
  assign _04263_ = _04262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6528" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1017];
  assign _04264_ = _04263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6528" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1018];
  assign _04265_ = _04264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6529" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1019];
  assign _04266_ = _04265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6529" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1020];
  assign _04267_ = _04266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6530" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva[1021];
  assign _04268_ = _04267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6530" *) _00856_;
  assign _04269_ = IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6536" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1];
  assign _04270_ = _04269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6536" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[2];
  assign _04271_ = _04270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6537" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[3];
  assign _04272_ = _04271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6537" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[4];
  assign _04273_ = _04272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6538" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[5];
  assign _04274_ = _04273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6538" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[6];
  assign _04275_ = _04274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6539" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[7];
  assign _04276_ = _04275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6539" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[8];
  assign _04277_ = _04276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6540" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[9];
  assign _04278_ = _04277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6540" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[10];
  assign _04279_ = _04278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6541" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[11];
  assign _04280_ = _04279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6541" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[12];
  assign _04281_ = _04280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6542" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[13];
  assign _04282_ = _04281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6542" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[14];
  assign _04283_ = _04282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6543" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[15];
  assign _04284_ = _04283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6543" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[16];
  assign _04285_ = _04284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6544" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[17];
  assign _04286_ = _04285_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6544" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[18];
  assign _04287_ = _04286_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6545" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[19];
  assign _04288_ = _04287_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6545" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[20];
  assign _04289_ = _04288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6546" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[21];
  assign _04290_ = _04289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6546" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[22];
  assign _04291_ = _04290_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6547" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[23];
  assign _04292_ = _04291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6547" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[24];
  assign _04293_ = _04292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6548" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[25];
  assign _04294_ = _04293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6548" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[26];
  assign _04295_ = _04294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6549" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[27];
  assign _04296_ = _04295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6549" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[28];
  assign _04297_ = _04296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6550" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[29];
  assign _04298_ = _04297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6550" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[30];
  assign _04299_ = _04298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6551" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[31];
  assign _04300_ = _04299_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6551" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[32];
  assign _04301_ = _04300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6552" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[33];
  assign _04302_ = _04301_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6552" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[34];
  assign _04303_ = _04302_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6553" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[35];
  assign _04304_ = _04303_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6553" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[36];
  assign _04305_ = _04304_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6554" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[37];
  assign _04306_ = _04305_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6554" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[38];
  assign _04307_ = _04306_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6555" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[39];
  assign _04308_ = _04307_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6555" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[40];
  assign _04309_ = _04308_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6556" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[41];
  assign _04310_ = _04309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6556" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[42];
  assign _04311_ = _04310_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6557" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[43];
  assign _04312_ = _04311_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6557" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[44];
  assign _04313_ = _04312_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6558" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[45];
  assign _04314_ = _04313_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6558" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[46];
  assign _04315_ = _04314_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6559" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[47];
  assign _04316_ = _04315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6559" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[48];
  assign _04317_ = _04316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6560" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[49];
  assign _04318_ = _04317_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6560" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[50];
  assign _04319_ = _04318_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6561" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[51];
  assign _04320_ = _04319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6561" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[52];
  assign _04321_ = _04320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6562" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[53];
  assign _04322_ = _04321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6562" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[54];
  assign _04323_ = _04322_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6563" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[55];
  assign _04324_ = _04323_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6563" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[56];
  assign _04325_ = _04324_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6564" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[57];
  assign _04326_ = _04325_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6564" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[58];
  assign _04327_ = _04326_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6565" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[59];
  assign _04328_ = _04327_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6565" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[60];
  assign _04329_ = _04328_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6566" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[61];
  assign _04330_ = _04329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6566" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[62];
  assign _04331_ = _04330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6567" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[63];
  assign _04332_ = _04331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6567" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[64];
  assign _04333_ = _04332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6568" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[65];
  assign _04334_ = _04333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6568" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[66];
  assign _04335_ = _04334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6569" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[67];
  assign _04336_ = _04335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6569" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[68];
  assign _04337_ = _04336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6570" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[69];
  assign _04338_ = _04337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6570" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[70];
  assign _04339_ = _04338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6571" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[71];
  assign _04340_ = _04339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6571" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[72];
  assign _04341_ = _04340_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6572" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[73];
  assign _04342_ = _04341_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6572" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[74];
  assign _04343_ = _04342_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6573" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[75];
  assign _04344_ = _04343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6573" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[76];
  assign _04345_ = _04344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6574" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[77];
  assign _04346_ = _04345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6574" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[78];
  assign _04347_ = _04346_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6575" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[79];
  assign _04348_ = _04347_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6575" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[80];
  assign _04349_ = _04348_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6576" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[81];
  assign _04350_ = _04349_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6576" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[82];
  assign _04351_ = _04350_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6577" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[83];
  assign _04352_ = _04351_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6577" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[84];
  assign _04353_ = _04352_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6578" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[85];
  assign _04354_ = _04353_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6578" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[86];
  assign _04355_ = _04354_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6579" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[87];
  assign _04356_ = _04355_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6579" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[88];
  assign _04357_ = _04356_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6580" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[89];
  assign _04358_ = _04357_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6580" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[90];
  assign _04359_ = _04358_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6581" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[91];
  assign _04360_ = _04359_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6581" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[92];
  assign _04361_ = _04360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6582" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[93];
  assign _04362_ = _04361_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6582" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[94];
  assign _04363_ = _04362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6583" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[95];
  assign _04364_ = _04363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6583" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[96];
  assign _04365_ = _04364_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6584" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[97];
  assign _04366_ = _04365_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6584" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[98];
  assign _04367_ = _04366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6585" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[99];
  assign _04368_ = _04367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6585" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[100];
  assign _04369_ = _04368_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6586" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[101];
  assign _04370_ = _04369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6586" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[102];
  assign _04371_ = _04370_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6587" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[103];
  assign _04372_ = _04371_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6587" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[104];
  assign _04373_ = _04372_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6588" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[105];
  assign _04374_ = _04373_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6588" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[106];
  assign _04375_ = _04374_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6589" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[107];
  assign _04376_ = _04375_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6589" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[108];
  assign _04377_ = _04376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6590" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[109];
  assign _04378_ = _04377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6590" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[110];
  assign _04379_ = _04378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6591" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[111];
  assign _04380_ = _04379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6591" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[112];
  assign _04381_ = _04380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6592" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[113];
  assign _04382_ = _04381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6592" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[114];
  assign _04383_ = _04382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6593" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[115];
  assign _04384_ = _04383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6593" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[116];
  assign _04385_ = _04384_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6594" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[117];
  assign _04386_ = _04385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6594" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[118];
  assign _04387_ = _04386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6595" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[119];
  assign _04388_ = _04387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6595" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[120];
  assign _04389_ = _04388_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6596" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[121];
  assign _04390_ = _04389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6596" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[122];
  assign _04391_ = _04390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6597" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[123];
  assign _04392_ = _04391_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6597" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[124];
  assign _04393_ = _04392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6598" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[125];
  assign _04394_ = _04393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6598" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[126];
  assign _04395_ = _04394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6599" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[127];
  assign _04396_ = _04395_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6599" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[128];
  assign _04397_ = _04396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6600" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[129];
  assign _04398_ = _04397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6600" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[130];
  assign _04399_ = _04398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6601" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[131];
  assign _04400_ = _04399_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6601" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[132];
  assign _04401_ = _04400_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6602" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[133];
  assign _04402_ = _04401_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6602" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[134];
  assign _04403_ = _04402_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6603" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[135];
  assign _04404_ = _04403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6603" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[136];
  assign _04405_ = _04404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6604" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[137];
  assign _04406_ = _04405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6604" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[138];
  assign _04407_ = _04406_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6605" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[139];
  assign _04408_ = _04407_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6605" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[140];
  assign _04409_ = _04408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6606" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[141];
  assign _04410_ = _04409_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6606" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[142];
  assign _04411_ = _04410_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6607" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[143];
  assign _04412_ = _04411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6607" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[144];
  assign _04413_ = _04412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6608" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[145];
  assign _04414_ = _04413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6608" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[146];
  assign _04415_ = _04414_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6609" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[147];
  assign _04416_ = _04415_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6609" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[148];
  assign _04417_ = _04416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6610" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[149];
  assign _04418_ = _04417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6610" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[150];
  assign _04419_ = _04418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6611" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[151];
  assign _04420_ = _04419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6611" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[152];
  assign _04421_ = _04420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6612" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[153];
  assign _04422_ = _04421_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6612" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[154];
  assign _04423_ = _04422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6613" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[155];
  assign _04424_ = _04423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6613" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[156];
  assign _04425_ = _04424_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6614" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[157];
  assign _04426_ = _04425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6614" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[158];
  assign _04427_ = _04426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6615" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[159];
  assign _04428_ = _04427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6615" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[160];
  assign _04429_ = _04428_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6616" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[161];
  assign _04430_ = _04429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6616" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[162];
  assign _04431_ = _04430_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6617" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[163];
  assign _04432_ = _04431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6617" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[164];
  assign _04433_ = _04432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6618" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[165];
  assign _04434_ = _04433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6618" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[166];
  assign _04435_ = _04434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6619" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[167];
  assign _04436_ = _04435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6619" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[168];
  assign _04437_ = _04436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6620" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[169];
  assign _04438_ = _04437_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6620" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[170];
  assign _04439_ = _04438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6621" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[171];
  assign _04440_ = _04439_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6621" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[172];
  assign _04441_ = _04440_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6622" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[173];
  assign _04442_ = _04441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6622" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[174];
  assign _04443_ = _04442_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6623" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[175];
  assign _04444_ = _04443_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6623" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[176];
  assign _04445_ = _04444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6624" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[177];
  assign _04446_ = _04445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6624" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[178];
  assign _04447_ = _04446_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6625" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[179];
  assign _04448_ = _04447_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6625" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[180];
  assign _04449_ = _04448_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6626" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[181];
  assign _04450_ = _04449_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6626" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[182];
  assign _04451_ = _04450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6627" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[183];
  assign _04452_ = _04451_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6627" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[184];
  assign _04453_ = _04452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6628" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[185];
  assign _04454_ = _04453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6628" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[186];
  assign _04455_ = _04454_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6629" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[187];
  assign _04456_ = _04455_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6629" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[188];
  assign _04457_ = _04456_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6630" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[189];
  assign _04458_ = _04457_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6630" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[190];
  assign _04459_ = _04458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6631" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[191];
  assign _04460_ = _04459_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6631" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[192];
  assign _04461_ = _04460_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6632" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[193];
  assign _04462_ = _04461_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6632" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[194];
  assign _04463_ = _04462_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6633" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[195];
  assign _04464_ = _04463_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6633" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[196];
  assign _04465_ = _04464_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6634" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[197];
  assign _04466_ = _04465_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6634" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[198];
  assign _04467_ = _04466_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6635" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[199];
  assign _04468_ = _04467_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6635" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[200];
  assign _04469_ = _04468_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6636" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[201];
  assign _04470_ = _04469_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6636" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[202];
  assign _04471_ = _04470_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6637" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[203];
  assign _04472_ = _04471_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6637" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[204];
  assign _04473_ = _04472_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6638" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[205];
  assign _04474_ = _04473_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6638" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[206];
  assign _04475_ = _04474_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6639" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[207];
  assign _04476_ = _04475_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6639" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[208];
  assign _04477_ = _04476_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6640" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[209];
  assign _04478_ = _04477_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6640" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[210];
  assign _04479_ = _04478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6641" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[211];
  assign _04480_ = _04479_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6641" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[212];
  assign _04481_ = _04480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6642" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[213];
  assign _04482_ = _04481_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6642" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[214];
  assign _04483_ = _04482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6643" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[215];
  assign _04484_ = _04483_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6643" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[216];
  assign _04485_ = _04484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6644" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[217];
  assign _04486_ = _04485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6644" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[218];
  assign _04487_ = _04486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6645" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[219];
  assign _04488_ = _04487_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6645" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[220];
  assign _04489_ = _04488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6646" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[221];
  assign _04490_ = _04489_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6646" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[222];
  assign _04491_ = _04490_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6647" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[223];
  assign _04492_ = _04491_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6647" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[224];
  assign _04493_ = _04492_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6648" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[225];
  assign _04494_ = _04493_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6648" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[226];
  assign _04495_ = _04494_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6649" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[227];
  assign _04496_ = _04495_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6649" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[228];
  assign _04497_ = _04496_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6650" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[229];
  assign _04498_ = _04497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6650" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[230];
  assign _04499_ = _04498_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6651" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[231];
  assign _04500_ = _04499_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6651" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[232];
  assign _04501_ = _04500_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6652" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[233];
  assign _04502_ = _04501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6652" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[234];
  assign _04503_ = _04502_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6653" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[235];
  assign _04504_ = _04503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6653" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[236];
  assign _04505_ = _04504_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6654" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[237];
  assign _04506_ = _04505_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6654" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[238];
  assign _04507_ = _04506_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6655" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[239];
  assign _04508_ = _04507_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6655" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[240];
  assign _04509_ = _04508_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6656" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[241];
  assign _04510_ = _04509_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6656" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[242];
  assign _04511_ = _04510_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6657" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[243];
  assign _04512_ = _04511_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6657" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[244];
  assign _04513_ = _04512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6658" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[245];
  assign _04514_ = _04513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6658" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[246];
  assign _04515_ = _04514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6659" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[247];
  assign _04516_ = _04515_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6659" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[248];
  assign _04517_ = _04516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6660" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[249];
  assign _04518_ = _04517_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6660" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[250];
  assign _04519_ = _04518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6661" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[251];
  assign _04520_ = _04519_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6661" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[252];
  assign _04521_ = _04520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6662" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[253];
  assign _04522_ = _04521_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6662" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[254];
  assign _04523_ = _04522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6663" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[255];
  assign _04524_ = _04523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6663" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[256];
  assign _04525_ = _04524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6664" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[257];
  assign _04526_ = _04525_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6664" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[258];
  assign _04527_ = _04526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6665" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[259];
  assign _04528_ = _04527_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6665" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[260];
  assign _04529_ = _04528_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6666" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[261];
  assign _04530_ = _04529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6666" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[262];
  assign _04531_ = _04530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6667" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[263];
  assign _04532_ = _04531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6667" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[264];
  assign _04533_ = _04532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6668" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[265];
  assign _04534_ = _04533_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6668" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[266];
  assign _04535_ = _04534_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6669" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[267];
  assign _04536_ = _04535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6669" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[268];
  assign _04537_ = _04536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6670" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[269];
  assign _04538_ = _04537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6670" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[270];
  assign _04539_ = _04538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6671" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[271];
  assign _04540_ = _04539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6671" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[272];
  assign _04541_ = _04540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6672" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[273];
  assign _04542_ = _04541_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6672" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[274];
  assign _04543_ = _04542_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6673" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[275];
  assign _04544_ = _04543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6673" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[276];
  assign _04545_ = _04544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6674" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[277];
  assign _04546_ = _04545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6674" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[278];
  assign _04547_ = _04546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6675" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[279];
  assign _04548_ = _04547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6675" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[280];
  assign _04549_ = _04548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6676" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[281];
  assign _04550_ = _04549_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6676" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[282];
  assign _04551_ = _04550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6677" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[283];
  assign _04552_ = _04551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6677" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[284];
  assign _04553_ = _04552_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6678" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[285];
  assign _04554_ = _04553_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6678" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[286];
  assign _04555_ = _04554_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6679" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[287];
  assign _04556_ = _04555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6679" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[288];
  assign _04557_ = _04556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6680" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[289];
  assign _04558_ = _04557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6680" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[290];
  assign _04559_ = _04558_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6681" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[291];
  assign _04560_ = _04559_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6681" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[292];
  assign _04561_ = _04560_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6682" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[293];
  assign _04562_ = _04561_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6682" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[294];
  assign _04563_ = _04562_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6683" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[295];
  assign _04564_ = _04563_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6683" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[296];
  assign _04565_ = _04564_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6684" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[297];
  assign _04566_ = _04565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6684" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[298];
  assign _04567_ = _04566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6685" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[299];
  assign _04568_ = _04567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6685" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[300];
  assign _04569_ = _04568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6686" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[301];
  assign _04570_ = _04569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6686" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[302];
  assign _04571_ = _04570_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6687" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[303];
  assign _04572_ = _04571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6687" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[304];
  assign _04573_ = _04572_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6688" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[305];
  assign _04574_ = _04573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6688" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[306];
  assign _04575_ = _04574_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6689" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[307];
  assign _04576_ = _04575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6689" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[308];
  assign _04577_ = _04576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6690" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[309];
  assign _04578_ = _04577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6690" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[310];
  assign _04579_ = _04578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6691" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[311];
  assign _04580_ = _04579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6691" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[312];
  assign _04581_ = _04580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6692" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[313];
  assign _04582_ = _04581_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6692" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[314];
  assign _04583_ = _04582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6693" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[315];
  assign _04584_ = _04583_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6693" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[316];
  assign _04585_ = _04584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6694" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[317];
  assign _04586_ = _04585_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6694" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[318];
  assign _04587_ = _04586_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6695" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[319];
  assign _04588_ = _04587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6695" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[320];
  assign _04589_ = _04588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6696" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[321];
  assign _04590_ = _04589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6696" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[322];
  assign _04591_ = _04590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6697" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[323];
  assign _04592_ = _04591_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6697" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[324];
  assign _04593_ = _04592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6698" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[325];
  assign _04594_ = _04593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6698" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[326];
  assign _04595_ = _04594_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6699" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[327];
  assign _04596_ = _04595_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6699" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[328];
  assign _04597_ = _04596_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6700" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[329];
  assign _04598_ = _04597_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6700" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[330];
  assign _04599_ = _04598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6701" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[331];
  assign _04600_ = _04599_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6701" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[332];
  assign _04601_ = _04600_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6702" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[333];
  assign _04602_ = _04601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6702" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[334];
  assign _04603_ = _04602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6703" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[335];
  assign _04604_ = _04603_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6703" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[336];
  assign _04605_ = _04604_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6704" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[337];
  assign _04606_ = _04605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6704" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[338];
  assign _04607_ = _04606_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6705" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[339];
  assign _04608_ = _04607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6705" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[340];
  assign _04609_ = _04608_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6706" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[341];
  assign _04610_ = _04609_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6706" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[342];
  assign _04611_ = _04610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6707" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[343];
  assign _04612_ = _04611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6707" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[344];
  assign _04613_ = _04612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6708" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[345];
  assign _04614_ = _04613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6708" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[346];
  assign _04615_ = _04614_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6709" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[347];
  assign _04616_ = _04615_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6709" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[348];
  assign _04617_ = _04616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6710" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[349];
  assign _04618_ = _04617_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6710" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[350];
  assign _04619_ = _04618_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6711" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[351];
  assign _04620_ = _04619_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6711" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[352];
  assign _04621_ = _04620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6712" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[353];
  assign _04622_ = _04621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6712" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[354];
  assign _04623_ = _04622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6713" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[355];
  assign _04624_ = _04623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6713" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[356];
  assign _04625_ = _04624_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6714" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[357];
  assign _04626_ = _04625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6714" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[358];
  assign _04627_ = _04626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6715" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[359];
  assign _04628_ = _04627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6715" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[360];
  assign _04629_ = _04628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6716" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[361];
  assign _04630_ = _04629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6716" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[362];
  assign _04631_ = _04630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6717" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[363];
  assign _04632_ = _04631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6717" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[364];
  assign _04633_ = _04632_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6718" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[365];
  assign _04634_ = _04633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6718" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[366];
  assign _04635_ = _04634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6719" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[367];
  assign _04636_ = _04635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6719" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[368];
  assign _04637_ = _04636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6720" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[369];
  assign _04638_ = _04637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6720" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[370];
  assign _04639_ = _04638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6721" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[371];
  assign _04640_ = _04639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6721" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[372];
  assign _04641_ = _04640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6722" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[373];
  assign _04642_ = _04641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6722" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[374];
  assign _04643_ = _04642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6723" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[375];
  assign _04644_ = _04643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6723" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[376];
  assign _04645_ = _04644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6724" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[377];
  assign _04646_ = _04645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6724" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[378];
  assign _04647_ = _04646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6725" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[379];
  assign _04648_ = _04647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6725" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[380];
  assign _04649_ = _04648_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6726" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[381];
  assign _04650_ = _04649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6726" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[382];
  assign _04651_ = _04650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6727" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[383];
  assign _04652_ = _04651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6727" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[384];
  assign _04653_ = _04652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6728" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[385];
  assign _04654_ = _04653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6728" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[386];
  assign _04655_ = _04654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6729" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[387];
  assign _04656_ = _04655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6729" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[388];
  assign _04657_ = _04656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6730" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[389];
  assign _04658_ = _04657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6730" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[390];
  assign _04659_ = _04658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6731" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[391];
  assign _04660_ = _04659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6731" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[392];
  assign _04661_ = _04660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6732" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[393];
  assign _04662_ = _04661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6732" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[394];
  assign _04663_ = _04662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6733" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[395];
  assign _04664_ = _04663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6733" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[396];
  assign _04665_ = _04664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6734" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[397];
  assign _04666_ = _04665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6734" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[398];
  assign _04667_ = _04666_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6735" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[399];
  assign _04668_ = _04667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6735" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[400];
  assign _04669_ = _04668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6736" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[401];
  assign _04670_ = _04669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6736" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[402];
  assign _04671_ = _04670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6737" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[403];
  assign _04672_ = _04671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6737" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[404];
  assign _04673_ = _04672_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6738" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[405];
  assign _04674_ = _04673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6738" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[406];
  assign _04675_ = _04674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6739" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[407];
  assign _04676_ = _04675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6739" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[408];
  assign _04677_ = _04676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6740" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[409];
  assign _04678_ = _04677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6740" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[410];
  assign _04679_ = _04678_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6741" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[411];
  assign _04680_ = _04679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6741" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[412];
  assign _04681_ = _04680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6742" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[413];
  assign _04682_ = _04681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6742" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[414];
  assign _04683_ = _04682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6743" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[415];
  assign _04684_ = _04683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6743" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[416];
  assign _04685_ = _04684_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6744" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[417];
  assign _04686_ = _04685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6744" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[418];
  assign _04687_ = _04686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6745" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[419];
  assign _04688_ = _04687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6745" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[420];
  assign _04689_ = _04688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6746" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[421];
  assign _04690_ = _04689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6746" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[422];
  assign _04691_ = _04690_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6747" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[423];
  assign _04692_ = _04691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6747" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[424];
  assign _04693_ = _04692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6748" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[425];
  assign _04694_ = _04693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6748" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[426];
  assign _04695_ = _04694_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6749" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[427];
  assign _04696_ = _04695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6749" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[428];
  assign _04697_ = _04696_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6750" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[429];
  assign _04698_ = _04697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6750" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[430];
  assign _04699_ = _04698_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6751" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[431];
  assign _04700_ = _04699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6751" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[432];
  assign _04701_ = _04700_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6752" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[433];
  assign _04702_ = _04701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6752" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[434];
  assign _04703_ = _04702_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6753" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[435];
  assign _04704_ = _04703_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6753" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[436];
  assign _04705_ = _04704_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6754" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[437];
  assign _04706_ = _04705_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6754" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[438];
  assign _04707_ = _04706_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6755" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[439];
  assign _04708_ = _04707_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6755" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[440];
  assign _04709_ = _04708_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6756" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[441];
  assign _04710_ = _04709_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6756" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[442];
  assign _04711_ = _04710_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6757" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[443];
  assign _04712_ = _04711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6757" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[444];
  assign _04713_ = _04712_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6758" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[445];
  assign _04714_ = _04713_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6758" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[446];
  assign _04715_ = _04714_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6759" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[447];
  assign _04716_ = _04715_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6759" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[448];
  assign _04717_ = _04716_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6760" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[449];
  assign _04718_ = _04717_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6760" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[450];
  assign _04719_ = _04718_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6761" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[451];
  assign _04720_ = _04719_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6761" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[452];
  assign _04721_ = _04720_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6762" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[453];
  assign _04722_ = _04721_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6762" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[454];
  assign _04723_ = _04722_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6763" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[455];
  assign _04724_ = _04723_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6763" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[456];
  assign _04725_ = _04724_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6764" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[457];
  assign _04726_ = _04725_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6764" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[458];
  assign _04727_ = _04726_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6765" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[459];
  assign _04728_ = _04727_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6765" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[460];
  assign _04729_ = _04728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6766" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[461];
  assign _04730_ = _04729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6766" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[462];
  assign _04731_ = _04730_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6767" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[463];
  assign _04732_ = _04731_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6767" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[464];
  assign _04733_ = _04732_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6768" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[465];
  assign _04734_ = _04733_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6768" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[466];
  assign _04735_ = _04734_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6769" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[467];
  assign _04736_ = _04735_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6769" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[468];
  assign _04737_ = _04736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6770" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[469];
  assign _04738_ = _04737_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6770" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[470];
  assign _04739_ = _04738_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6771" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[471];
  assign _04740_ = _04739_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6771" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[472];
  assign _04741_ = _04740_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6772" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[473];
  assign _04742_ = _04741_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6772" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[474];
  assign _04743_ = _04742_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6773" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[475];
  assign _04744_ = _04743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6773" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[476];
  assign _04745_ = _04744_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6774" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[477];
  assign _04746_ = _04745_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6774" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[478];
  assign _04747_ = _04746_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6775" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[479];
  assign _04748_ = _04747_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6775" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[480];
  assign _04749_ = _04748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6776" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[481];
  assign _04750_ = _04749_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6776" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[482];
  assign _04751_ = _04750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6777" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[483];
  assign _04752_ = _04751_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6777" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[484];
  assign _04753_ = _04752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6778" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[485];
  assign _04754_ = _04753_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6778" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[486];
  assign _04755_ = _04754_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6779" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[487];
  assign _04756_ = _04755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6779" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[488];
  assign _04757_ = _04756_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6780" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[489];
  assign _04758_ = _04757_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6780" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[490];
  assign _04759_ = _04758_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6781" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[491];
  assign _04760_ = _04759_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6781" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[492];
  assign _04761_ = _04760_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6782" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[493];
  assign _04762_ = _04761_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6782" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[494];
  assign _04763_ = _04762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6783" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[495];
  assign _04764_ = _04763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6783" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[496];
  assign _04765_ = _04764_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6784" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[497];
  assign _04766_ = _04765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6784" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[498];
  assign _04767_ = _04766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6785" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[499];
  assign _04768_ = _04767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6785" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[500];
  assign _04769_ = _04768_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6786" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[501];
  assign _04770_ = _04769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6786" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[502];
  assign _04771_ = _04770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6787" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[503];
  assign _04772_ = _04771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6787" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[504];
  assign _04773_ = _04772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6788" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[505];
  assign _04774_ = _04773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6788" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[506];
  assign _04775_ = _04774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6789" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[507];
  assign _04776_ = _04775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6789" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[508];
  assign _04777_ = _04776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6790" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[509];
  assign _04778_ = _04777_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6790" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[510];
  assign _04779_ = _04778_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6791" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[511];
  assign _04780_ = _04779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6791" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[512];
  assign _04781_ = _04780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6792" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[513];
  assign _04782_ = _04781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6792" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[514];
  assign _04783_ = _04782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6793" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[515];
  assign _04784_ = _04783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6793" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[516];
  assign _04785_ = _04784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6794" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[517];
  assign _04786_ = _04785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6794" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[518];
  assign _04787_ = _04786_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6795" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[519];
  assign _04788_ = _04787_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6795" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[520];
  assign _04789_ = _04788_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6796" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[521];
  assign _04790_ = _04789_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6796" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[522];
  assign _04791_ = _04790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6797" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[523];
  assign _04792_ = _04791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6797" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[524];
  assign _04793_ = _04792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6798" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[525];
  assign _04794_ = _04793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6798" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[526];
  assign _04795_ = _04794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6799" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[527];
  assign _04796_ = _04795_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6799" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[528];
  assign _04797_ = _04796_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6800" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[529];
  assign _04798_ = _04797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6800" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[530];
  assign _04799_ = _04798_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6801" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[531];
  assign _04800_ = _04799_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6801" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[532];
  assign _04801_ = _04800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6802" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[533];
  assign _04802_ = _04801_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6802" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[534];
  assign _04803_ = _04802_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6803" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[535];
  assign _04804_ = _04803_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6803" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[536];
  assign _04805_ = _04804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6804" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[537];
  assign _04806_ = _04805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6804" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[538];
  assign _04807_ = _04806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6805" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[539];
  assign _04808_ = _04807_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6805" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[540];
  assign _04809_ = _04808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6806" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[541];
  assign _04810_ = _04809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6806" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[542];
  assign _04811_ = _04810_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6807" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[543];
  assign _04812_ = _04811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6807" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[544];
  assign _04813_ = _04812_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6808" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[545];
  assign _04814_ = _04813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6808" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[546];
  assign _04815_ = _04814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6809" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[547];
  assign _04816_ = _04815_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6809" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[548];
  assign _04817_ = _04816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6810" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[549];
  assign _04818_ = _04817_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6810" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[550];
  assign _04819_ = _04818_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6811" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[551];
  assign _04820_ = _04819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6811" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[552];
  assign _04821_ = _04820_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6812" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[553];
  assign _04822_ = _04821_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6812" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[554];
  assign _04823_ = _04822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6813" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[555];
  assign _04824_ = _04823_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6813" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[556];
  assign _04825_ = _04824_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6814" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[557];
  assign _04826_ = _04825_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6814" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[558];
  assign _04827_ = _04826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6815" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[559];
  assign _04828_ = _04827_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6815" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[560];
  assign _04829_ = _04828_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6816" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[561];
  assign _04830_ = _04829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6816" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[562];
  assign _04831_ = _04830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6817" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[563];
  assign _04832_ = _04831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6817" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[564];
  assign _04833_ = _04832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6818" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[565];
  assign _04834_ = _04833_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6818" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[566];
  assign _04835_ = _04834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6819" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[567];
  assign _04836_ = _04835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6819" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[568];
  assign _04837_ = _04836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6820" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[569];
  assign _04838_ = _04837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6820" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[570];
  assign _04839_ = _04838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6821" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[571];
  assign _04840_ = _04839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6821" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[572];
  assign _04841_ = _04840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6822" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[573];
  assign _04842_ = _04841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6822" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[574];
  assign _04843_ = _04842_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6823" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[575];
  assign _04844_ = _04843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6823" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[576];
  assign _04845_ = _04844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6824" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[577];
  assign _04846_ = _04845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6824" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[578];
  assign _04847_ = _04846_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6825" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[579];
  assign _04848_ = _04847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6825" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[580];
  assign _04849_ = _04848_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6826" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[581];
  assign _04850_ = _04849_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6826" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[582];
  assign _04851_ = _04850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6827" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[583];
  assign _04852_ = _04851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6827" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[584];
  assign _04853_ = _04852_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6828" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[585];
  assign _04854_ = _04853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6828" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[586];
  assign _04855_ = _04854_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6829" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[587];
  assign _04856_ = _04855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6829" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[588];
  assign _04857_ = _04856_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6830" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[589];
  assign _04858_ = _04857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6830" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[590];
  assign _04859_ = _04858_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6831" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[591];
  assign _04860_ = _04859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6831" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[592];
  assign _04861_ = _04860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6832" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[593];
  assign _04862_ = _04861_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6832" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[594];
  assign _04863_ = _04862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6833" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[595];
  assign _04864_ = _04863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6833" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[596];
  assign _04865_ = _04864_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6834" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[597];
  assign _04866_ = _04865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6834" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[598];
  assign _04867_ = _04866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6835" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[599];
  assign _04868_ = _04867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6835" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[600];
  assign _04869_ = _04868_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6836" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[601];
  assign _04870_ = _04869_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6836" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[602];
  assign _04871_ = _04870_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6837" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[603];
  assign _04872_ = _04871_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6837" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[604];
  assign _04873_ = _04872_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6838" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[605];
  assign _04874_ = _04873_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6838" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[606];
  assign _04875_ = _04874_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6839" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[607];
  assign _04876_ = _04875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6839" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[608];
  assign _04877_ = _04876_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6840" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[609];
  assign _04878_ = _04877_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6840" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[610];
  assign _04879_ = _04878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6841" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[611];
  assign _04880_ = _04879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6841" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[612];
  assign _04881_ = _04880_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6842" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[613];
  assign _04882_ = _04881_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6842" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[614];
  assign _04883_ = _04882_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6843" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[615];
  assign _04884_ = _04883_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6843" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[616];
  assign _04885_ = _04884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6844" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[617];
  assign _04886_ = _04885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6844" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[618];
  assign _04887_ = _04886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6845" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[619];
  assign _04888_ = _04887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6845" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[620];
  assign _04889_ = _04888_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6846" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[621];
  assign _04890_ = _04889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6846" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[622];
  assign _04891_ = _04890_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6847" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[623];
  assign _04892_ = _04891_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6847" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[624];
  assign _04893_ = _04892_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6848" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[625];
  assign _04894_ = _04893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6848" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[626];
  assign _04895_ = _04894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6849" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[627];
  assign _04896_ = _04895_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6849" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[628];
  assign _04897_ = _04896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6850" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[629];
  assign _04898_ = _04897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6850" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[630];
  assign _04899_ = _04898_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6851" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[631];
  assign _04900_ = _04899_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6851" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[632];
  assign _04901_ = _04900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6852" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[633];
  assign _04902_ = _04901_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6852" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[634];
  assign _04903_ = _04902_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6853" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[635];
  assign _04904_ = _04903_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6853" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[636];
  assign _04905_ = _04904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6854" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[637];
  assign _04906_ = _04905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6854" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[638];
  assign _04907_ = _04906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6855" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[639];
  assign _04908_ = _04907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6855" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[640];
  assign _04909_ = _04908_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6856" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[641];
  assign _04910_ = _04909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6856" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[642];
  assign _04911_ = _04910_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6857" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[643];
  assign _04912_ = _04911_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6857" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[644];
  assign _04913_ = _04912_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6858" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[645];
  assign _04914_ = _04913_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6858" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[646];
  assign _04915_ = _04914_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6859" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[647];
  assign _04916_ = _04915_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6859" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[648];
  assign _04917_ = _04916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6860" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[649];
  assign _04918_ = _04917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6860" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[650];
  assign _04919_ = _04918_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6861" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[651];
  assign _04920_ = _04919_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6861" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[652];
  assign _04921_ = _04920_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6862" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[653];
  assign _04922_ = _04921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6862" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[654];
  assign _04923_ = _04922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6863" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[655];
  assign _04924_ = _04923_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6863" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[656];
  assign _04925_ = _04924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6864" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[657];
  assign _04926_ = _04925_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6864" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[658];
  assign _04927_ = _04926_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6865" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[659];
  assign _04928_ = _04927_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6865" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[660];
  assign _04929_ = _04928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6866" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[661];
  assign _04930_ = _04929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6866" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[662];
  assign _04931_ = _04930_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6867" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[663];
  assign _04932_ = _04931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6867" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[664];
  assign _04933_ = _04932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6868" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[665];
  assign _04934_ = _04933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6868" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[666];
  assign _04935_ = _04934_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6869" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[667];
  assign _04936_ = _04935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6869" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[668];
  assign _04937_ = _04936_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6870" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[669];
  assign _04938_ = _04937_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6870" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[670];
  assign _04939_ = _04938_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6871" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[671];
  assign _04940_ = _04939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6871" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[672];
  assign _04941_ = _04940_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6872" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[673];
  assign _04942_ = _04941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6872" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[674];
  assign _04943_ = _04942_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6873" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[675];
  assign _04944_ = _04943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6873" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[676];
  assign _04945_ = _04944_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6874" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[677];
  assign _04946_ = _04945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6874" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[678];
  assign _04947_ = _04946_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6875" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[679];
  assign _04948_ = _04947_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6875" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[680];
  assign _04949_ = _04948_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6876" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[681];
  assign _04950_ = _04949_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6876" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[682];
  assign _04951_ = _04950_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6877" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[683];
  assign _04952_ = _04951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6877" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[684];
  assign _04953_ = _04952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6878" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[685];
  assign _04954_ = _04953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6878" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[686];
  assign _04955_ = _04954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6879" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[687];
  assign _04956_ = _04955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6879" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[688];
  assign _04957_ = _04956_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6880" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[689];
  assign _04958_ = _04957_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6880" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[690];
  assign _04959_ = _04958_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6881" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[691];
  assign _04960_ = _04959_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6881" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[692];
  assign _04961_ = _04960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6882" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[693];
  assign _04962_ = _04961_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6882" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[694];
  assign _04963_ = _04962_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6883" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[695];
  assign _04964_ = _04963_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6883" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[696];
  assign _04965_ = _04964_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6884" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[697];
  assign _04966_ = _04965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6884" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[698];
  assign _04967_ = _04966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6885" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[699];
  assign _04968_ = _04967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6885" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[700];
  assign _04969_ = _04968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6886" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[701];
  assign _04970_ = _04969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6886" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[702];
  assign _04971_ = _04970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6887" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[703];
  assign _04972_ = _04971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6887" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[704];
  assign _04973_ = _04972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6888" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[705];
  assign _04974_ = _04973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6888" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[706];
  assign _04975_ = _04974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6889" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[707];
  assign _04976_ = _04975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6889" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[708];
  assign _04977_ = _04976_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6890" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[709];
  assign _04978_ = _04977_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6890" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[710];
  assign _04979_ = _04978_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6891" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[711];
  assign _04980_ = _04979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6891" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[712];
  assign _04981_ = _04980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6892" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[713];
  assign _04982_ = _04981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6892" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[714];
  assign _04983_ = _04982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6893" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[715];
  assign _04984_ = _04983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6893" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[716];
  assign _04985_ = _04984_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6894" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[717];
  assign _04986_ = _04985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6894" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[718];
  assign _04987_ = _04986_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6895" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[719];
  assign _04988_ = _04987_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6895" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[720];
  assign _04989_ = _04988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6896" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[721];
  assign _04990_ = _04989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6896" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[722];
  assign _04991_ = _04990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6897" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[723];
  assign _04992_ = _04991_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6897" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[724];
  assign _04993_ = _04992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6898" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[725];
  assign _04994_ = _04993_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6898" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[726];
  assign _04995_ = _04994_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6899" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[727];
  assign _04996_ = _04995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6899" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[728];
  assign _04997_ = _04996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6900" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[729];
  assign _04998_ = _04997_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6900" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[730];
  assign _04999_ = _04998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6901" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[731];
  assign _05000_ = _04999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6901" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[732];
  assign _05001_ = _05000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6902" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[733];
  assign _05002_ = _05001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6902" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[734];
  assign _05003_ = _05002_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6903" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[735];
  assign _05004_ = _05003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6903" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[736];
  assign _05005_ = _05004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6904" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[737];
  assign _05006_ = _05005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6904" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[738];
  assign _05007_ = _05006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6905" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[739];
  assign _05008_ = _05007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6905" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[740];
  assign _05009_ = _05008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6906" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[741];
  assign _05010_ = _05009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6906" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[742];
  assign _05011_ = _05010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6907" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[743];
  assign _05012_ = _05011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6907" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[744];
  assign _05013_ = _05012_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6908" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[745];
  assign _05014_ = _05013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6908" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[746];
  assign _05015_ = _05014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6909" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[747];
  assign _05016_ = _05015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6909" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[748];
  assign _05017_ = _05016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6910" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[749];
  assign _05018_ = _05017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6910" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[750];
  assign _05019_ = _05018_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6911" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[751];
  assign _05020_ = _05019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6911" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[752];
  assign _05021_ = _05020_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6912" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[753];
  assign _05022_ = _05021_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6912" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[754];
  assign _05023_ = _05022_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6913" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[755];
  assign _05024_ = _05023_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6913" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[756];
  assign _05025_ = _05024_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6914" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[757];
  assign _05026_ = _05025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6914" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[758];
  assign _05027_ = _05026_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6915" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[759];
  assign _05028_ = _05027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6915" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[760];
  assign _05029_ = _05028_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6916" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[761];
  assign _05030_ = _05029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6916" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[762];
  assign _05031_ = _05030_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6917" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[763];
  assign _05032_ = _05031_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6917" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[764];
  assign _05033_ = _05032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6918" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[765];
  assign _05034_ = _05033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6918" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[766];
  assign _05035_ = _05034_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6919" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[767];
  assign _05036_ = _05035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6919" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[768];
  assign _05037_ = _05036_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6920" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[769];
  assign _05038_ = _05037_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6920" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[770];
  assign _05039_ = _05038_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6921" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[771];
  assign _05040_ = _05039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6921" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[772];
  assign _05041_ = _05040_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6922" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[773];
  assign _05042_ = _05041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6922" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[774];
  assign _05043_ = _05042_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6923" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[775];
  assign _05044_ = _05043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6923" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[776];
  assign _05045_ = _05044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6924" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[777];
  assign _05046_ = _05045_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6924" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[778];
  assign _05047_ = _05046_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6925" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[779];
  assign _05048_ = _05047_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6925" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[780];
  assign _05049_ = _05048_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6926" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[781];
  assign _05050_ = _05049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6926" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[782];
  assign _05051_ = _05050_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6927" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[783];
  assign _05052_ = _05051_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6927" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[784];
  assign _05053_ = _05052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6928" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[785];
  assign _05054_ = _05053_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6928" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[786];
  assign _05055_ = _05054_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6929" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[787];
  assign _05056_ = _05055_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6929" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[788];
  assign _05057_ = _05056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6930" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[789];
  assign _05058_ = _05057_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6930" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[790];
  assign _05059_ = _05058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6931" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[791];
  assign _05060_ = _05059_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6931" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[792];
  assign _05061_ = _05060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6932" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[793];
  assign _05062_ = _05061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6932" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[794];
  assign _05063_ = _05062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6933" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[795];
  assign _05064_ = _05063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6933" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[796];
  assign _05065_ = _05064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6934" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[797];
  assign _05066_ = _05065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6934" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[798];
  assign _05067_ = _05066_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6935" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[799];
  assign _05068_ = _05067_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6935" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[800];
  assign _05069_ = _05068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6936" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[801];
  assign _05070_ = _05069_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6936" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[802];
  assign _05071_ = _05070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6937" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[803];
  assign _05072_ = _05071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6937" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[804];
  assign _05073_ = _05072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6938" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[805];
  assign _05074_ = _05073_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6938" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[806];
  assign _05075_ = _05074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6939" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[807];
  assign _05076_ = _05075_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6939" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[808];
  assign _05077_ = _05076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6940" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[809];
  assign _05078_ = _05077_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6940" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[810];
  assign _05079_ = _05078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6941" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[811];
  assign _05080_ = _05079_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6941" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[812];
  assign _05081_ = _05080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6942" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[813];
  assign _05082_ = _05081_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6942" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[814];
  assign _05083_ = _05082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6943" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[815];
  assign _05084_ = _05083_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6943" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[816];
  assign _05085_ = _05084_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6944" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[817];
  assign _05086_ = _05085_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6944" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[818];
  assign _05087_ = _05086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6945" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[819];
  assign _05088_ = _05087_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6945" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[820];
  assign _05089_ = _05088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6946" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[821];
  assign _05090_ = _05089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6946" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[822];
  assign _05091_ = _05090_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6947" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[823];
  assign _05092_ = _05091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6947" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[824];
  assign _05093_ = _05092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6948" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[825];
  assign _05094_ = _05093_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6948" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[826];
  assign _05095_ = _05094_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6949" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[827];
  assign _05096_ = _05095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6949" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[828];
  assign _05097_ = _05096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6950" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[829];
  assign _05098_ = _05097_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6950" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[830];
  assign _05099_ = _05098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6951" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[831];
  assign _05100_ = _05099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6951" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[832];
  assign _05101_ = _05100_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6952" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[833];
  assign _05102_ = _05101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6952" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[834];
  assign _05103_ = _05102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6953" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[835];
  assign _05104_ = _05103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6953" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[836];
  assign _05105_ = _05104_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6954" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[837];
  assign _05106_ = _05105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6954" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[838];
  assign _05107_ = _05106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6955" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[839];
  assign _05108_ = _05107_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6955" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[840];
  assign _05109_ = _05108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6956" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[841];
  assign _05110_ = _05109_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6956" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[842];
  assign _05111_ = _05110_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6957" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[843];
  assign _05112_ = _05111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6957" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[844];
  assign _05113_ = _05112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6958" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[845];
  assign _05114_ = _05113_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6958" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[846];
  assign _05115_ = _05114_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6959" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[847];
  assign _05116_ = _05115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6959" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[848];
  assign _05117_ = _05116_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6960" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[849];
  assign _05118_ = _05117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6960" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[850];
  assign _05119_ = _05118_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6961" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[851];
  assign _05120_ = _05119_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6961" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[852];
  assign _05121_ = _05120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6962" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[853];
  assign _05122_ = _05121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6962" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[854];
  assign _05123_ = _05122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6963" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[855];
  assign _05124_ = _05123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6963" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[856];
  assign _05125_ = _05124_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6964" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[857];
  assign _05126_ = _05125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6964" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[858];
  assign _05127_ = _05126_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6965" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[859];
  assign _05128_ = _05127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6965" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[860];
  assign _05129_ = _05128_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6966" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[861];
  assign _05130_ = _05129_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6966" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[862];
  assign _05131_ = _05130_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6967" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[863];
  assign _05132_ = _05131_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6967" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[864];
  assign _05133_ = _05132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6968" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[865];
  assign _05134_ = _05133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6968" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[866];
  assign _05135_ = _05134_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6969" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[867];
  assign _05136_ = _05135_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6969" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[868];
  assign _05137_ = _05136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6970" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[869];
  assign _05138_ = _05137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6970" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[870];
  assign _05139_ = _05138_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6971" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[871];
  assign _05140_ = _05139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6971" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[872];
  assign _05141_ = _05140_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6972" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[873];
  assign _05142_ = _05141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6972" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[874];
  assign _05143_ = _05142_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6973" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[875];
  assign _05144_ = _05143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6973" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[876];
  assign _05145_ = _05144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6974" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[877];
  assign _05146_ = _05145_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6974" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[878];
  assign _05147_ = _05146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6975" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[879];
  assign _05148_ = _05147_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6975" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[880];
  assign _05149_ = _05148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6976" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[881];
  assign _05150_ = _05149_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6976" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[882];
  assign _05151_ = _05150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6977" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[883];
  assign _05152_ = _05151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6977" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[884];
  assign _05153_ = _05152_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6978" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[885];
  assign _05154_ = _05153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6978" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[886];
  assign _05155_ = _05154_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6979" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[887];
  assign _05156_ = _05155_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6979" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[888];
  assign _05157_ = _05156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6980" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[889];
  assign _05158_ = _05157_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6980" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[890];
  assign _05159_ = _05158_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6981" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[891];
  assign _05160_ = _05159_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6981" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[892];
  assign _05161_ = _05160_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6982" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[893];
  assign _05162_ = _05161_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6982" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[894];
  assign _05163_ = _05162_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6983" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[895];
  assign _05164_ = _05163_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6983" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[896];
  assign _05165_ = _05164_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6984" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[897];
  assign _05166_ = _05165_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6984" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[898];
  assign _05167_ = _05166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6985" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[899];
  assign _05168_ = _05167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6985" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[900];
  assign _05169_ = _05168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6986" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[901];
  assign _05170_ = _05169_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6986" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[902];
  assign _05171_ = _05170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6987" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[903];
  assign _05172_ = _05171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6987" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[904];
  assign _05173_ = _05172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6988" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[905];
  assign _05174_ = _05173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6988" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[906];
  assign _05175_ = _05174_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6989" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[907];
  assign _05176_ = _05175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6989" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[908];
  assign _05177_ = _05176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6990" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[909];
  assign _05178_ = _05177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6990" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[910];
  assign _05179_ = _05178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6991" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[911];
  assign _05180_ = _05179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6991" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[912];
  assign _05181_ = _05180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6992" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[913];
  assign _05182_ = _05181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6992" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[914];
  assign _05183_ = _05182_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6993" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[915];
  assign _05184_ = _05183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6993" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[916];
  assign _05185_ = _05184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6994" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[917];
  assign _05186_ = _05185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6994" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[918];
  assign _05187_ = _05186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6995" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[919];
  assign _05188_ = _05187_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6995" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[920];
  assign _05189_ = _05188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6996" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[921];
  assign _05190_ = _05189_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6996" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[922];
  assign _05191_ = _05190_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6997" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[923];
  assign _05192_ = _05191_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6997" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[924];
  assign _05193_ = _05192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6998" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[925];
  assign _05194_ = _05193_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6998" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[926];
  assign _05195_ = _05194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6999" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[927];
  assign _05196_ = _05195_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:6999" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[928];
  assign _05197_ = _05196_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7000" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[929];
  assign _05198_ = _05197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7000" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[930];
  assign _05199_ = _05198_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7001" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[931];
  assign _05200_ = _05199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7001" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[932];
  assign _05201_ = _05200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7002" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[933];
  assign _05202_ = _05201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7002" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[934];
  assign _05203_ = _05202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7003" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[935];
  assign _05204_ = _05203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7003" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[936];
  assign _05205_ = _05204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7004" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[937];
  assign _05206_ = _05205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7004" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[938];
  assign _05207_ = _05206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7005" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[939];
  assign _05208_ = _05207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7005" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[940];
  assign _05209_ = _05208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7006" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[941];
  assign _05210_ = _05209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7006" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[942];
  assign _05211_ = _05210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7007" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[943];
  assign _05212_ = _05211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7007" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[944];
  assign _05213_ = _05212_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7008" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[945];
  assign _05214_ = _05213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7008" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[946];
  assign _05215_ = _05214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7009" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[947];
  assign _05216_ = _05215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7009" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[948];
  assign _05217_ = _05216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7010" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[949];
  assign _05218_ = _05217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7010" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[950];
  assign _05219_ = _05218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7011" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[951];
  assign _05220_ = _05219_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7011" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[952];
  assign _05221_ = _05220_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7012" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[953];
  assign _05222_ = _05221_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7012" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[954];
  assign _05223_ = _05222_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7013" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[955];
  assign _05224_ = _05223_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7013" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[956];
  assign _05225_ = _05224_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7014" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[957];
  assign _05226_ = _05225_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7014" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[958];
  assign _05227_ = _05226_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7015" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[959];
  assign _05228_ = _05227_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7015" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[960];
  assign _05229_ = _05228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7016" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[961];
  assign _05230_ = _05229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7016" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[962];
  assign _05231_ = _05230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7017" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[963];
  assign _05232_ = _05231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7017" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[964];
  assign _05233_ = _05232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7018" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[965];
  assign _05234_ = _05233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7018" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[966];
  assign _05235_ = _05234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7019" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[967];
  assign _05236_ = _05235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7019" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[968];
  assign _05237_ = _05236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7020" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[969];
  assign _05238_ = _05237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7020" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[970];
  assign _05239_ = _05238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7021" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[971];
  assign _05240_ = _05239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7021" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[972];
  assign _05241_ = _05240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7022" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[973];
  assign _05242_ = _05241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7022" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[974];
  assign _05243_ = _05242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7023" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[975];
  assign _05244_ = _05243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7023" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[976];
  assign _05245_ = _05244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7024" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[977];
  assign _05246_ = _05245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7024" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[978];
  assign _05247_ = _05246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7025" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[979];
  assign _05248_ = _05247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7025" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[980];
  assign _05249_ = _05248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7026" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[981];
  assign _05250_ = _05249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7026" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[982];
  assign _05251_ = _05250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7027" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[983];
  assign _05252_ = _05251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7027" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[984];
  assign _05253_ = _05252_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7028" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[985];
  assign _05254_ = _05253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7028" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[986];
  assign _05255_ = _05254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7029" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[987];
  assign _05256_ = _05255_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7029" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[988];
  assign _05257_ = _05256_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7030" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[989];
  assign _05258_ = _05257_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7030" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[990];
  assign _05259_ = _05258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7031" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[991];
  assign _05260_ = _05259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7031" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[992];
  assign _05261_ = _05260_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7032" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[993];
  assign _05262_ = _05261_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7032" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[994];
  assign _05263_ = _05262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7033" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[995];
  assign _05264_ = _05263_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7033" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[996];
  assign _05265_ = _05264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7034" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[997];
  assign _05266_ = _05265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7034" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[998];
  assign _05267_ = _05266_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7035" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[999];
  assign _05268_ = _05267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7035" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1000];
  assign _05269_ = _05268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7036" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1001];
  assign _05270_ = _05269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7036" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1002];
  assign _05271_ = _05270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7037" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1003];
  assign _05272_ = _05271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7037" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1004];
  assign _05273_ = _05272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7038" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1005];
  assign _05274_ = _05273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7038" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1006];
  assign _05275_ = _05274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7039" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1007];
  assign _05276_ = _05275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7039" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1008];
  assign _05277_ = _05276_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7040" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1009];
  assign _05278_ = _05277_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7040" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1010];
  assign _05279_ = _05278_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7041" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1011];
  assign _05280_ = _05279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7041" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1012];
  assign _05281_ = _05280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7042" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1013];
  assign _05282_ = _05281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7042" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1014];
  assign _05283_ = _05282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7043" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1015];
  assign _05284_ = _05283_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7043" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1016];
  assign _05285_ = _05284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7044" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1017];
  assign _05286_ = _05285_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7044" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1018];
  assign _05287_ = _05286_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7045" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1019];
  assign _05288_ = _05287_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7045" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1020];
  assign _05289_ = _05288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7046" *) IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva[1021];
  assign _05290_ = _05289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7046" *) _00857_;
  assign asn_158 = mul_mul_land_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7090" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign asn_162 = mul_mul_land_1_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7093" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign asn_166 = mul_mul_land_3_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7096" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign asn_170 = mul_mul_land_2_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7099" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign or_tmp_1 = io_read_cfg_mul_bypass_rsc_svs_st_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7110" *) mul_mul_land_1_lpi_1_dfm_st_1;
  assign _05291_ = mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl[9] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7112" *) IsZero_8U_23U_land_1_lpi_1_dfm_4;
  assign _05292_ = _05291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7112" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp;
  assign or_19_nl = _05292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7112" *) _00862_;
  assign _05293_ = or_tmp_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7114" *) mux_5_nl;
  assign or_tmp_59 = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7116" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign _05294_ = or_tmp_59 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7116" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  assign _05295_ = _05294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7117" *) _00768_;
  assign _05296_ = _05295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7117" *) _00766_;
  assign _05297_ = _05296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7117" *) _00765_;
  assign _05298_ = _05297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7117" *) chn_mul_out_rsci_bawt;
  assign _05299_ = mul_mul_land_1_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7120" *) _00765_;
  assign _05300_ = _05299_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7120" *) chn_mul_out_rsci_bawt;
  assign _05301_ = _05300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7120" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign or_26_nl = _05301_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7120" *) _00766_;
  assign _05302_ = or_tmp_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7123" *) IsZero_8U_23U_land_1_lpi_1_dfm_4;
  assign _05303_ = _05302_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7124" *) mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign or_tmp_12 = _05303_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7124" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp;
  assign or_tmp_15 = io_read_cfg_mul_bypass_rsc_svs_st_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7125" *) mul_mul_land_2_lpi_1_dfm_st_1;
  assign _05304_ = mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl[9] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7127" *) IsZero_8U_23U_land_2_lpi_1_dfm_4;
  assign _05305_ = _05304_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7127" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp;
  assign or_34_nl = _05305_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7127" *) _00863_;
  assign _05306_ = or_tmp_15 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7129" *) mux_10_nl;
  assign or_tmp_75 = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7131" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign _05307_ = or_tmp_75 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7131" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  assign _05308_ = _05307_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7132" *) _00772_;
  assign _05309_ = _05308_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7132" *) _00766_;
  assign _05310_ = _05309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7132" *) _00765_;
  assign _05311_ = _05310_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7132" *) chn_mul_out_rsci_bawt;
  assign _05312_ = mul_mul_land_2_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7135" *) _00765_;
  assign _05313_ = _05312_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7135" *) chn_mul_out_rsci_bawt;
  assign _05314_ = _05313_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7135" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign or_40_nl = _05314_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7135" *) _00766_;
  assign _05315_ = or_tmp_15 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7138" *) IsZero_8U_23U_land_2_lpi_1_dfm_4;
  assign _05316_ = _05315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7139" *) mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign or_tmp_26 = _05316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7139" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp;
  assign or_tmp_29 = io_read_cfg_mul_bypass_rsc_svs_st_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7140" *) mul_mul_land_3_lpi_1_dfm_st_1;
  assign _05317_ = mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl[9] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7142" *) IsZero_8U_23U_land_3_lpi_1_dfm_4;
  assign _05318_ = _05317_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7142" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp;
  assign or_48_nl = _05318_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7142" *) _00864_;
  assign _05319_ = or_tmp_29 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7144" *) mux_15_nl;
  assign or_tmp_91 = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7146" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign _05320_ = or_tmp_91 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7146" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  assign _05321_ = _05320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7147" *) _00776_;
  assign _05322_ = _05321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7147" *) _00766_;
  assign _05323_ = _05322_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7147" *) _00765_;
  assign _05324_ = _05323_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7147" *) chn_mul_out_rsci_bawt;
  assign _05325_ = mul_mul_land_3_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7150" *) _00765_;
  assign _05326_ = _05325_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7150" *) chn_mul_out_rsci_bawt;
  assign _05327_ = _05326_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7150" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign or_54_nl = _05327_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7150" *) _00766_;
  assign _05328_ = or_tmp_29 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7153" *) IsZero_8U_23U_land_3_lpi_1_dfm_4;
  assign _05329_ = _05328_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7154" *) mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign or_tmp_40 = _05329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7154" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp;
  assign _05330_ = mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl[9] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7156" *) IsZero_8U_23U_land_lpi_1_dfm_4;
  assign _05331_ = _05330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7156" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp;
  assign _05332_ = _05331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7157" *) _00865_;
  assign _05333_ = _05332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7157" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05334_ = _05333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7157" *) mul_mul_land_lpi_1_dfm_st_1;
  assign or_498_nl = _00866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7159" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st;
  assign _05335_ = or_498_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7159" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05336_ = _05335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7159" *) mul_mul_land_lpi_1_dfm_st_1;
  assign or_tmp_107 = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7162" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05337_ = or_tmp_107 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7162" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign _05338_ = _05337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7163" *) _00780_;
  assign _05339_ = _05338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7163" *) _00766_;
  assign _05340_ = _05339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7163" *) _00765_;
  assign _05341_ = _05340_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7163" *) chn_mul_out_rsci_bawt;
  assign or_tmp_46 = mul_mul_land_lpi_1_dfm_st_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7165" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05342_ = or_74_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7167" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05343_ = _05342_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7167" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign or_65_nl = _05343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7167" *) _00766_;
  assign _05344_ = or_tmp_46 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7170" *) mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign _05345_ = _05344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7171" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp;
  assign or_tmp_51 = _05345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7171" *) IsZero_8U_23U_land_lpi_1_dfm_4;
  assign _05346_ = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7177" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign or_tmp_123 = _05346_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7177" *) mul_mul_land_1_lpi_1_dfm_5;
  assign or_tmp_128 = FpMul_8U_23U_FpMul_8U_23U_and_itm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7178" *) FpMul_8U_23U_lor_6_lpi_1_dfm_6;
  assign or_tmp_132 = _00458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7181" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2;
  assign _05347_ = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7184" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _05348_ = _05347_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7184" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign or_tmp_146 = _05348_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7184" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05349_ = nor_143_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7185" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign or_tmp_167 = _05349_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7185" *) _00766_;
  assign or_189_cse = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7187" *) _00766_;
  assign _05350_ = mul_mul_land_1_lpi_1_dfm_st_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7190" *) _00765_;
  assign _05351_ = _05350_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7190" *) chn_mul_out_rsci_bawt;
  assign _05352_ = _05351_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7190" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign or_187_nl = _05352_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7190" *) _00752_;
  assign or_193_nl = mul_mul_land_1_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7194" *) mul_mul_land_1_lpi_1_dfm_st_5;
  assign _05353_ = or_193_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7194" *) _00765_;
  assign _05354_ = _05353_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7194" *) chn_mul_out_rsci_bawt;
  assign _05355_ = _05354_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7195" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _05356_ = _05355_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7195" *) _00752_;
  assign _05357_ = nor_143_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7196" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05358_ = _05357_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7197" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05359_ = _05358_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7197" *) _00766_;
  assign _05360_ = mul_mul_land_1_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7199" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05361_ = _05360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7199" *) _00766_;
  assign _05362_ = or_tmp_59 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7206" *) _00766_;
  assign _05363_ = _05362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7206" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _05364_ = _05363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7207" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign _05365_ = _05364_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7207" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05366_ = _01027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7209" *) IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  assign _05367_ = _05366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7209" *) mul_mul_land_1_lpi_1_dfm_st_5;
  assign _05368_ = _05367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7209" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign _05369_ = or_744_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7212" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05370_ = _05369_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7212" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign or_tmp_211 = _05370_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7212" *) mul_mul_land_2_lpi_1_dfm_5;
  assign or_tmp_216 = FpMul_8U_23U_FpMul_8U_23U_and_12_itm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7213" *) FpMul_8U_23U_lor_7_lpi_1_dfm_6;
  assign _05371_ = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7215" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _05372_ = _05371_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7215" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign or_tmp_235 = _05372_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7215" *) mul_mul_land_2_lpi_1_dfm_5;
  assign or_tmp_252 = FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7216" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign _05373_ = mul_mul_land_2_lpi_1_dfm_st_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7218" *) _00765_;
  assign _05374_ = _05373_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7218" *) chn_mul_out_rsci_bawt;
  assign _05375_ = _05374_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7218" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign or_tmp_256 = _05375_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7218" *) _00752_;
  assign _05376_ = _05374_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7221" *) mul_mul_land_2_lpi_1_dfm_6;
  assign _05377_ = _05376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7222" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _05378_ = _05377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7222" *) _00752_;
  assign _05379_ = nor_143_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7223" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05380_ = _05379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7224" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05381_ = _05380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7224" *) _00766_;
  assign _05382_ = mul_mul_land_2_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7226" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05383_ = _05382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7226" *) _00766_;
  assign _05384_ = asn_170 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7228" *) _00752_;
  assign _05385_ = or_tmp_75 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7233" *) _00766_;
  assign _05386_ = _05385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7233" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _05387_ = _05386_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7234" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign _05388_ = _05387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7234" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05389_ = _01031_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7236" *) IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  assign _05390_ = _05389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7236" *) mul_mul_land_2_lpi_1_dfm_st_5;
  assign _05391_ = _05390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7236" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _05392_ = or_745_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7240" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05393_ = _05392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7240" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign or_tmp_291 = _05393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7240" *) mul_mul_land_3_lpi_1_dfm_5;
  assign or_tmp_296 = FpMul_8U_23U_FpMul_8U_23U_and_13_itm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7241" *) FpMul_8U_23U_lor_8_lpi_1_dfm_6;
  assign _05394_ = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7243" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _05395_ = _05394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7243" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign or_tmp_315 = _05395_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7243" *) mul_mul_land_3_lpi_1_dfm_5;
  assign or_tmp_332 = FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7244" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign _05396_ = mul_mul_land_3_lpi_1_dfm_st_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7246" *) _00765_;
  assign _05397_ = _05396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7246" *) chn_mul_out_rsci_bawt;
  assign _05398_ = _05397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7246" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign or_tmp_336 = _05398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7246" *) _00752_;
  assign _05399_ = _05397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7249" *) mul_mul_land_3_lpi_1_dfm_6;
  assign _05400_ = _05399_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7250" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _05401_ = _05400_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7250" *) _00752_;
  assign _05402_ = nor_143_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7251" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05403_ = _05402_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7252" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05404_ = _05403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7252" *) _00766_;
  assign _05405_ = mul_mul_land_3_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7254" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05406_ = _05405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7254" *) _00766_;
  assign _05407_ = asn_166 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7256" *) _00752_;
  assign _05408_ = or_tmp_91 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7261" *) _00766_;
  assign _05409_ = _05408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7261" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _05410_ = _05409_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7262" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign _05411_ = _05410_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7262" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05412_ = _01035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7264" *) IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  assign _05413_ = _05412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7264" *) mul_mul_land_3_lpi_1_dfm_st_5;
  assign _05414_ = _05413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7264" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign _05415_ = or_430_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7268" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05416_ = _05415_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7268" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign or_tmp_371 = _05416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7268" *) mul_mul_land_lpi_1_dfm_5;
  assign or_tmp_376 = FpMul_8U_23U_FpMul_8U_23U_and_14_itm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7269" *) FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  assign _05417_ = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7273" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _05418_ = _05417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7273" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign or_tmp_395 = _05418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7273" *) mul_mul_land_lpi_1_dfm_5;
  assign _05419_ = nor_143_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7274" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05420_ = _05419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7275" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign or_tmp_411 = _05420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7275" *) _00766_;
  assign _05421_ = mul_mul_land_lpi_1_dfm_st_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7277" *) _00765_;
  assign _05422_ = _05421_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7277" *) chn_mul_out_rsci_bawt;
  assign _05423_ = _05422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7277" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign or_tmp_415 = _05423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7277" *) _00752_;
  assign or_435_nl = or_tmp_107 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7278" *) _00766_;
  assign _05424_ = nor_143_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7281" *) mul_mul_land_lpi_1_dfm_5;
  assign _05425_ = _05424_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7282" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05426_ = _05425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7282" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05427_ = _05426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7282" *) _00766_;
  assign _05428_ = mul_mul_land_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7284" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05429_ = _05428_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7284" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05430_ = _05429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7284" *) _00766_;
  assign _05431_ = asn_158 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7286" *) _00752_;
  assign _05432_ = or_435_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7290" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _05433_ = _05432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7291" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign _05434_ = _05433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7291" *) mul_mul_land_lpi_1_dfm_5;
  assign _05435_ = _01039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7293" *) IsNaN_8U_23U_land_lpi_1_dfm_8;
  assign _05436_ = _05435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7293" *) mul_mul_land_lpi_1_dfm_st_5;
  assign _05437_ = _05436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7293" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _05438_ = chn_mul_in_rsci_d_mxwt[95] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7296" *) chn_mul_in_rsci_d_mxwt[31];
  assign _05439_ = _05438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7296" *) chn_mul_in_rsci_d_mxwt[63];
  assign _05440_ = _05439_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7296" *) chn_mul_in_rsci_d_mxwt[127];
  assign _05441_ = _05440_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7296" *) _00828_;
  assign or_tmp_461 = _00867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7297" *) cfg_mul_bypass_rsci_d;
  assign or_tmp_517 = FpMul_8U_23U_FpMul_8U_23U_and_14_itm | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7304" *) _00868_;
  assign or_dcpl_8 = cfg_mul_bypass_rsci_d | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7311" *) _00784_;
  assign or_dcpl_13 = and_dcpl_23 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7314" *) _00766_;
  assign _05442_ = or_dcpl_13 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7337" *) or_tmp_59;
  assign _05443_ = _05442_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7338" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  assign _05444_ = _05443_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7339" *) _00768_;
  assign or_dcpl_22 = _05444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7339" *) or_27_cse;
  assign or_dcpl_23 = mul_mul_land_1_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7340" *) cfg_precision[0];
  assign or_dcpl_26 = or_189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7341" *) and_dcpl_23;
  assign _05445_ = or_dcpl_26 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7342" *) or_dcpl_23;
  assign or_dcpl_27 = _05445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7342" *) _00875_;
  assign _05446_ = or_dcpl_13 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7343" *) or_tmp_75;
  assign _05447_ = _05446_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7344" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  assign _05448_ = _05447_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7345" *) _00772_;
  assign or_dcpl_37 = _05448_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7345" *) or_27_cse;
  assign _05449_ = or_dcpl_26 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7346" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign or_dcpl_40 = _05449_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7346" *) or_27_cse;
  assign _05450_ = or_dcpl_13 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7347" *) or_tmp_91;
  assign _05451_ = _05450_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7348" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  assign _05452_ = _05451_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7349" *) _00776_;
  assign or_dcpl_50 = _05452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7349" *) or_27_cse;
  assign _05453_ = or_dcpl_26 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7350" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign or_dcpl_53 = _05453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7350" *) or_27_cse;
  assign _05454_ = or_189_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7351" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05455_ = _05454_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7351" *) and_dcpl_23;
  assign _05456_ = _05455_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7352" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign _05457_ = _05456_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7353" *) _00780_;
  assign or_dcpl_63 = _05457_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7353" *) or_27_cse;
  assign _05458_ = or_dcpl_26 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7354" *) mul_mul_land_lpi_1_dfm_st_4;
  assign or_dcpl_66 = _05458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7354" *) or_27_cse;
  assign _05459_ = or_tmp_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7360" *) cfg_precision[0];
  assign or_dcpl_99 = _05459_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7360" *) or_dcpl_96;
  assign _05460_ = or_tmp_15 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7361" *) cfg_precision[0];
  assign or_dcpl_102 = _05460_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7361" *) or_dcpl_96;
  assign _05461_ = or_tmp_29 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7362" *) cfg_precision[0];
  assign or_dcpl_105 = _05461_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7362" *) or_dcpl_96;
  assign _05462_ = or_tmp_46 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7363" *) cfg_precision[0];
  assign or_dcpl_108 = _05462_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7363" *) or_dcpl_96;
  assign or_dcpl_110 = _00784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7364" *) or_27_cse;
  assign or_dcpl_125 = and_dcpl_37 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7365" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign chn_mul_in_rsci_ld_core_psct_mx0c0 = and_20_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7369" *) fsm_output[0];
  assign _05463_ = or_dcpl_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7370" *) _00876_;
  assign _05464_ = and_dcpl_24 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7473" *) and_dcpl_26;
  assign _05465_ = or_tmp_588 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7481" *) chn_mul_op_rsci_ld_core_psct_mx0c1;
  assign _05466_ = or_tmp_591 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7489" *) main_stage_v_2_mx0c1;
  assign _05467_ = _00465_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7745" *) main_stage_v_3_mx0c1;
  assign _05468_ = or_tmp_587 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8382" *) main_stage_v_1_mx0c1;
  assign _05469_ = or_tmp_461 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8430" *) cfg_mul_src_rsci_d;
  assign _05470_ = _00530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8497" *) cfg_mul_src_1_sva_st_1_mx0c1;
  assign _05471_ = or_dcpl_27 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8539" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  assign _05472_ = _05449_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8605" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  assign _05473_ = _05472_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8605" *) or_27_cse;
  assign _05474_ = _05453_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8670" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  assign _05475_ = _05474_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8670" *) or_27_cse;
  assign _05476_ = _05458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8735" *) IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  assign _05477_ = _05476_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8735" *) or_27_cse;
  assign _05478_ = mul_mul_land_1_lpi_1_dfm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8776" *) mul_mul_land_1_lpi_1_dfm_st_1;
  assign _05479_ = _05478_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8776" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05480_ = and_135_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8784" *) mul_mul_if_and_6_rgt;
  assign _05481_ = _05480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8784" *) mul_mul_if_and_7_rgt;
  assign _05482_ = mul_mul_land_2_lpi_1_dfm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8804" *) mul_mul_land_2_lpi_1_dfm_st_1;
  assign _05483_ = _05482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8804" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05484_ = and_137_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8812" *) mul_mul_if_and_4_rgt;
  assign _05485_ = _05484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8812" *) mul_mul_if_and_5_rgt;
  assign _05486_ = mul_mul_land_3_lpi_1_dfm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8832" *) mul_mul_land_3_lpi_1_dfm_st_1;
  assign _05487_ = _05486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8832" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05488_ = and_139_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8840" *) mul_mul_if_and_2_rgt;
  assign _05489_ = _05488_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8840" *) mul_mul_if_and_3_rgt;
  assign _05490_ = mul_mul_land_lpi_1_dfm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8860" *) mul_mul_land_lpi_1_dfm_st_1;
  assign _05491_ = _05490_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8860" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05492_ = and_141_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8868" *) mul_mul_if_and_rgt;
  assign _05493_ = _05492_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8868" *) mul_mul_if_and_1_rgt;
  assign _05494_ = or_dcpl_26 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8879" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign _05495_ = _05494_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8880" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  assign _05496_ = _05495_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8880" *) or_27_cse;
  assign _05497_ = _00566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8890" *) and_146_rgt;
  assign _05498_ = _00571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8902" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05499_ = or_dcpl_26 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8911" *) or_tmp_252;
  assign _05500_ = _05499_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8911" *) or_27_cse;
  assign _05501_ = _00575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8921" *) and_150_rgt;
  assign _05502_ = or_dcpl_26 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8932" *) or_tmp_332;
  assign _05503_ = _05502_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8932" *) or_27_cse;
  assign _05504_ = _00580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8942" *) and_154_rgt;
  assign _05505_ = _05458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8954" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign _05506_ = _05505_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8954" *) or_27_cse;
  assign _05507_ = _00585_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8964" *) and_158_rgt;
  assign _05508_ = or_dcpl_99 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8983" *) fsm_output[0];
  assign _05509_ = or_dcpl_102 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8999" *) fsm_output[0];
  assign _05510_ = or_dcpl_105 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9015" *) fsm_output[0];
  assign _05511_ = or_dcpl_108 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9031" *) fsm_output[0];
  assign _05512_ = or_dcpl_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9079" *) fsm_output[0];
  assign _05513_ = FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05514_ = _05513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *) mul_mul_land_1_lpi_1_dfm_st_1;
  assign _05515_ = _05514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *) cfg_precision[0];
  assign _05516_ = _05515_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *) or_dcpl_96;
  assign _05517_ = _05516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9088" *) fsm_output[0];
  assign _05518_ = or_dcpl_125 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9097" *) mul_mul_land_1_lpi_1_dfm_st_1;
  assign _05519_ = _05518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9098" *) _00812_;
  assign _05520_ = _05519_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9098" *) fsm_output[0];
  assign _05521_ = FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05522_ = _05521_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *) mul_mul_land_2_lpi_1_dfm_st_1;
  assign _05523_ = _05522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *) cfg_precision[0];
  assign _05524_ = _05523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *) or_dcpl_96;
  assign _05525_ = _05524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9107" *) fsm_output[0];
  assign _05526_ = or_dcpl_125 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9116" *) mul_mul_land_2_lpi_1_dfm_st_1;
  assign _05527_ = _05526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9117" *) _00812_;
  assign _05528_ = _05527_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9117" *) fsm_output[0];
  assign _05529_ = FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05530_ = _05529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *) mul_mul_land_3_lpi_1_dfm_st_1;
  assign _05531_ = _05530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *) cfg_precision[0];
  assign _05532_ = _05531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *) or_dcpl_96;
  assign _05533_ = _05532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9126" *) fsm_output[0];
  assign _05534_ = or_dcpl_125 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9135" *) mul_mul_land_3_lpi_1_dfm_st_1;
  assign _05535_ = _05534_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9136" *) _00812_;
  assign _05536_ = _05535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9136" *) fsm_output[0];
  assign _05537_ = _01071_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9145" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05538_ = _05537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9145" *) mul_mul_land_lpi_1_dfm_st_1;
  assign _05539_ = _05538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9146" *) cfg_precision[0];
  assign _05540_ = _05539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9146" *) or_dcpl_96;
  assign _05541_ = _05540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9146" *) fsm_output[0];
  assign _05542_ = or_dcpl_125 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9154" *) mul_mul_land_lpi_1_dfm_st_1;
  assign _05543_ = _05542_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9155" *) _00812_;
  assign _05544_ = _05543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9155" *) fsm_output[0];
  assign _05545_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9161" *) IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_1_sva;
  assign _05546_ = _00929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9161" *) IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva;
  assign _05547_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9169" *) IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva;
  assign _05548_ = _00930_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9169" *) IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_1_sva;
  assign _05549_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9176" *) IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_2_sva;
  assign _05550_ = _00931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9176" *) IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva;
  assign _05551_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9184" *) IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva;
  assign _05552_ = _00932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9184" *) IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_2_sva;
  assign _05553_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9191" *) IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_3_sva;
  assign _05554_ = _00933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9191" *) IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva;
  assign _05555_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9199" *) IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva;
  assign _05556_ = _00934_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9199" *) IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_3_sva;
  assign _05557_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9205" *) IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_sva;
  assign _05558_ = _00935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9206" *) IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva;
  assign _05559_ = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1[31] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9213" *) IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva;
  assign _05560_ = _00936_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9214" *) IntShiftRight_64U_10U_32U_obits_fixed_nor_ovfl_sva;
  assign _05561_ = _01201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9224" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign or_839_nl = _00610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9236" *) asn_162;
  assign _05562_ = _01200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9242" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign or_838_nl = _00612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9254" *) asn_170;
  assign _05563_ = _01199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9260" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign or_837_nl = _00614_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9272" *) asn_166;
  assign _05564_ = _01198_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9278" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign or_836_nl = _00616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9290" *) asn_158;
  assign _05565_ = FpMul_8U_23U_lor_6_lpi_1_dfm_st | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9292" *) mul_mul_land_1_lpi_1_dfm_st_1;
  assign or_28_nl = _05565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9292" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05566_ = FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9295" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign _05567_ = _05566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9295" *) _00765_;
  assign _05568_ = _05567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9295" *) chn_mul_out_rsci_bawt;
  assign _05569_ = _05568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9296" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign or_31_nl = _05569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9296" *) _00766_;
  assign _05570_ = FpMul_8U_23U_lor_7_lpi_1_dfm_st | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9299" *) mul_mul_land_2_lpi_1_dfm_st_1;
  assign or_42_nl = _05570_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9299" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05571_ = or_tmp_252 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9302" *) _00765_;
  assign _05572_ = _05571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9302" *) chn_mul_out_rsci_bawt;
  assign _05573_ = _05572_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9303" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign or_45_nl = _05573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9303" *) _00766_;
  assign _05574_ = FpMul_8U_23U_lor_8_lpi_1_dfm_st | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9306" *) mul_mul_land_3_lpi_1_dfm_st_1;
  assign or_56_nl = _05574_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9306" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05575_ = or_tmp_332 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9309" *) _00765_;
  assign _05576_ = _05575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9309" *) chn_mul_out_rsci_bawt;
  assign _05577_ = _05576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9310" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign or_59_nl = _05577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9310" *) _00766_;
  assign _05578_ = FpMul_8U_23U_lor_1_lpi_1_dfm_st | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9313" *) mul_mul_land_lpi_1_dfm_st_1;
  assign or_67_nl = _05578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9313" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05579_ = FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9316" *) _00765_;
  assign _05580_ = _05579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9316" *) chn_mul_out_rsci_bawt;
  assign _05581_ = _05580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9316" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05582_ = _05581_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9317" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign or_70_nl = _05582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9317" *) _00766_;
  assign _05583_ = IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9320" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05584_ = _05583_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9320" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign _05585_ = _05584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9320" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05586_ = nor_301_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9321" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05587_ = _05586_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9322" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign or_142_nl = _05587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9322" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05588_ = _00941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9324" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05589_ = _05588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9324" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign or_143_nl = _05589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9324" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05590_ = _00942_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9327" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05591_ = _05590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9328" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign or_147_nl = _05591_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9328" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05592_ = _00617_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9331" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm;
  assign or_831_nl = _00943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9332" *) mux_37_nl;
  assign _05593_ = or_743_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9335" *) mux_38_nl;
  assign _05594_ = _01202_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9340" *) _00945_;
  assign or_153_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9343" *) _00946_;
  assign _05595_ = _05367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9347" *) mux_41_nl;
  assign _05596_ = _00767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9350" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05597_ = _05596_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9350" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign _05598_ = _05597_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9350" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  assign _05599_ = _05598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9350" *) nand_48_cse;
  assign _05600_ = _00947_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9352" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05601_ = _05600_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9352" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign _05602_ = _05601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9353" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  assign _05603_ = _05602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9353" *) nand_48_cse;
  assign _05604_ = or_tmp_173 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9356" *) mul_mul_land_1_lpi_1_dfm_st_5;
  assign _05605_ = _05604_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9356" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st_4;
  assign _05606_ = _05605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9357" *) _00948_;
  assign _05607_ = nor_301_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9359" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _05608_ = _05607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9360" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign or_165_nl = _05608_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9360" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05609_ = _00941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9362" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _05610_ = _05609_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9362" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign or_166_nl = _05610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9362" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05611_ = _00942_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9365" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _05612_ = _05611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9366" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign or_169_nl = _05612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9366" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05613_ = _05296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9371" *) mux_48_nl;
  assign _05614_ = _05368_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9374" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st_4;
  assign _05615_ = mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9375" *) FpMul_8U_23U_FpMul_8U_23U_nor_4_nl;
  assign _05616_ = _05614_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9375" *) _00949_;
  assign _05617_ = _05294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9378" *) nand_48_cse;
  assign _05618_ = _05605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9380" *) _00950_;
  assign _05619_ = FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9383" *) mul_mul_land_1_lpi_1_dfm_st_5;
  assign _05620_ = _05619_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9383" *) _00765_;
  assign _05621_ = _05620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9383" *) chn_mul_out_rsci_bawt;
  assign _05622_ = _05621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9384" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign or_181_nl = _05622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9384" *) _00752_;
  assign or_185_nl = mul_mul_land_1_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9385" *) or_tmp_167;
  assign _05623_ = nor_277_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9388" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign _05624_ = _05623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9388" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05625_ = FpMul_8U_23U_p_mant_p1_1_sva[47] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9390" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign _05626_ = _05625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9390" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05627_ = _00951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9395" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign or_210_nl = _05627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9395" *) mul_mul_land_1_lpi_1_dfm_5;
  assign or_211_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9397" *) mux_61_nl;
  assign _05628_ = _05362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9400" *) mux_62_nl;
  assign _05629_ = nor_282_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *) FpMul_8U_23U_lor_6_lpi_1_dfm_7;
  assign _05630_ = _05629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *) _00952_;
  assign _05631_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *) _00953_;
  assign _05632_ = _05367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9403" *) _00954_;
  assign _05633_ = nor_277_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9405" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05634_ = _05633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9406" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign _05635_ = _05634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9406" *) _00766_;
  assign _05636_ = _05635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9406" *) FpMul_8U_23U_lor_6_lpi_1_dfm_6;
  assign _05637_ = _05636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9407" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _05638_ = _05637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9407" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign _05639_ = _05638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9407" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05640_ = FpMul_8U_23U_p_mant_p1_1_sva[47] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9409" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05641_ = _05640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9409" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign _05642_ = _05641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9409" *) _00766_;
  assign _05643_ = _05642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9410" *) FpMul_8U_23U_lor_6_lpi_1_dfm_6;
  assign _05644_ = _05643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9410" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _05645_ = _05644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9410" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign _05646_ = _05645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9410" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05647_ = _00951_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9415" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05648_ = _05647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9415" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign _05649_ = _05648_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9415" *) _00766_;
  assign _05650_ = _05649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9416" *) FpMul_8U_23U_lor_6_lpi_1_dfm_6;
  assign _05651_ = _05650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9416" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _05652_ = _05651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9416" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign _05653_ = _05652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9416" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05654_ = nor_282_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9418" *) _00752_;
  assign _05655_ = _05654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9419" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _05656_ = _05655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9419" *) mul_mul_land_1_lpi_1_dfm_6;
  assign _05657_ = _05656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9419" *) IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  assign _05658_ = _05657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9420" *) mul_mul_land_1_lpi_1_dfm_st_5;
  assign _05659_ = _05658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9420" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign _05660_ = _05659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9420" *) FpMul_8U_23U_lor_6_lpi_1_dfm_7;
  assign _05661_ = _05660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9420" *) _00952_;
  assign _05662_ = IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9423" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign or_227_nl = _05662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9423" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05663_ = nor_264_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9424" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  assign _05664_ = _05663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9425" *) _00772_;
  assign _05665_ = _05664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9425" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign or_230_nl = _05665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9425" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05666_ = _00955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9427" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  assign _05667_ = _05666_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9428" *) _00772_;
  assign _05668_ = _05667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9428" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign or_231_nl = _05668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9428" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05669_ = _00956_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9431" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  assign _05670_ = _05669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9432" *) _00772_;
  assign _05671_ = _05670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9432" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign or_235_nl = _05671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9432" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05672_ = _00622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9435" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm;
  assign or_830_nl = _00957_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9436" *) mux_69_nl;
  assign _05673_ = _05385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9440" *) mux_71_nl;
  assign _05674_ = FpMul_8U_23U_lor_7_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9441" *) _00958_;
  assign _05675_ = nor_267_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9446" *) mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2;
  assign _05676_ = _05390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9451" *) mux_73_nl;
  assign _05677_ = _00771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9454" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05678_ = _05677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9454" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign _05679_ = _05678_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9454" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  assign _05680_ = _05679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9454" *) nand_45_cse;
  assign _05681_ = _00960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9456" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05682_ = _05681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9456" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign _05683_ = _05682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9457" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  assign _05684_ = _05683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9457" *) nand_45_cse;
  assign _05685_ = or_tmp_173 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9460" *) mul_mul_land_2_lpi_1_dfm_st_5;
  assign _05686_ = _05685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9460" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_4;
  assign _05687_ = _05686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9461" *) _00961_;
  assign _05688_ = nor_264_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9463" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _05689_ = _05688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9464" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign or_254_nl = _05689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9464" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05690_ = _00955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9466" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _05691_ = _05690_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9466" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign or_255_nl = _05691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9466" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05692_ = _00956_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9469" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _05693_ = _05692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9470" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign or_258_nl = _05693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9470" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05694_ = _05309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9475" *) mux_80_nl;
  assign _05695_ = _00962_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9477" *) _00752_;
  assign _05696_ = _05695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9477" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _05697_ = _05696_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9478" *) mul_mul_land_2_lpi_1_dfm_6;
  assign _05698_ = _05697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9478" *) IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  assign _05699_ = _05698_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9478" *) mul_mul_land_2_lpi_1_dfm_st_5;
  assign _05700_ = _05699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9479" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _05701_ = _05700_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9479" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_4;
  assign _05702_ = _05701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9479" *) _00958_;
  assign _05703_ = _05307_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9482" *) nand_45_cse;
  assign _05704_ = _05686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9484" *) _00958_;
  assign or_270_nl = or_tmp_252 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9486" *) or_tmp_167;
  assign _05705_ = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9490" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign _05706_ = _05705_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9490" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05707_ = nor_241_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9491" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05708_ = _05707_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9492" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign _05709_ = _05708_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9492" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05710_ = FpMul_8U_23U_p_mant_p1_2_sva[47] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9494" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05711_ = _05710_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9494" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign _05712_ = _05711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9494" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05713_ = _00963_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9499" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05714_ = _05713_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9499" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign or_292_nl = _05714_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9499" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05715_ = FpMul_8U_23U_lor_7_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9501" *) mux_91_nl;
  assign _05716_ = nor_245_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9507" *) FpMul_8U_23U_lor_7_lpi_1_dfm_7;
  assign _05717_ = _05716_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9507" *) _00965_;
  assign _05718_ = _00966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9508" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _05719_ = _05390_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9508" *) _00967_;
  assign _05720_ = _05707_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9511" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign _05721_ = _05720_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9511" *) _00766_;
  assign _05722_ = _05721_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9511" *) FpMul_8U_23U_lor_7_lpi_1_dfm_6;
  assign _05723_ = _05722_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9512" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _05724_ = _05723_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9512" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign _05725_ = _05724_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9512" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05726_ = _05710_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9514" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign _05727_ = _05726_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9514" *) _00766_;
  assign _05728_ = _05727_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9515" *) FpMul_8U_23U_lor_7_lpi_1_dfm_6;
  assign _05729_ = _05728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9515" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _05730_ = _05729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9515" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign _05731_ = _05730_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9515" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05732_ = _05713_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9520" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign _05733_ = _05732_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9520" *) _00766_;
  assign _05734_ = _05733_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9521" *) FpMul_8U_23U_lor_7_lpi_1_dfm_6;
  assign _05735_ = _05734_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9521" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _05736_ = _05735_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9521" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign _05737_ = _05736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9521" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05738_ = nor_245_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9523" *) _00752_;
  assign _05739_ = _05738_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9524" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _05740_ = _05739_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9524" *) mul_mul_land_2_lpi_1_dfm_6;
  assign _05741_ = _05740_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9524" *) IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  assign _05742_ = _05741_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9525" *) mul_mul_land_2_lpi_1_dfm_st_5;
  assign _05743_ = _05742_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9525" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _05744_ = _05743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9525" *) FpMul_8U_23U_lor_7_lpi_1_dfm_7;
  assign _05745_ = _05744_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9525" *) _00965_;
  assign _05746_ = IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9528" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign or_307_nl = _05746_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9528" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05747_ = nor_227_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9529" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  assign _05748_ = _05747_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9530" *) _00776_;
  assign _05749_ = _05748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9530" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign or_310_nl = _05749_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9530" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05750_ = _00968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9532" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  assign _05751_ = _05750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9533" *) _00776_;
  assign _05752_ = _05751_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9533" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign or_311_nl = _05752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9533" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05753_ = _00969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9536" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  assign _05754_ = _05753_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9537" *) _00776_;
  assign _05755_ = _05754_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9537" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign or_315_nl = _05755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9537" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05756_ = _00628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9540" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm;
  assign or_829_nl = _00970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9541" *) mux_100_nl;
  assign _05757_ = _05408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9545" *) mux_102_nl;
  assign _05758_ = FpMul_8U_23U_lor_8_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9546" *) _00971_;
  assign _05759_ = nor_230_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9551" *) mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2;
  assign _05760_ = _05413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9556" *) mux_104_nl;
  assign _05761_ = _00775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9559" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05762_ = _05761_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9559" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign _05763_ = _05762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9559" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  assign _05764_ = _05763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9559" *) nand_42_cse;
  assign _05765_ = _00973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9561" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05766_ = _05765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9561" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign _05767_ = _05766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9562" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  assign _05768_ = _05767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9562" *) nand_42_cse;
  assign _05769_ = or_tmp_173 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9565" *) mul_mul_land_3_lpi_1_dfm_st_5;
  assign _05770_ = _05769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9565" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_4;
  assign _05771_ = _05770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9566" *) _00974_;
  assign _05772_ = nor_227_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9568" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _05773_ = _05772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9569" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign or_334_nl = _05773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9569" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05774_ = _00968_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9571" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _05775_ = _05774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9571" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign or_335_nl = _05775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9571" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05776_ = _00969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9574" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _05777_ = _05776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9575" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign or_338_nl = _05777_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9575" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05778_ = _05322_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9580" *) mux_111_nl;
  assign _05779_ = _00975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9582" *) _00752_;
  assign _05780_ = _05779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9582" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _05781_ = _05780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9583" *) mul_mul_land_3_lpi_1_dfm_6;
  assign _05782_ = _05781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9583" *) IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  assign _05783_ = _05782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9583" *) mul_mul_land_3_lpi_1_dfm_st_5;
  assign _05784_ = _05783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9584" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign _05785_ = _05784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9584" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_4;
  assign _05786_ = _05785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9584" *) _00971_;
  assign _05787_ = _05320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9587" *) nand_42_cse;
  assign _05788_ = _05770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9589" *) _00971_;
  assign or_350_nl = or_tmp_332 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9591" *) or_tmp_167;
  assign _05789_ = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9595" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign _05790_ = _05789_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9595" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05791_ = nor_204_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9596" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05792_ = _05791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9597" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign _05793_ = _05792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9597" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05794_ = FpMul_8U_23U_p_mant_p1_3_sva[47] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9599" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05795_ = _05794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9599" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign _05796_ = _05795_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9599" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05797_ = _00976_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9604" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05798_ = _05797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9604" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign or_372_nl = _05798_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9604" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05799_ = FpMul_8U_23U_lor_8_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9606" *) mux_122_nl;
  assign _05800_ = nor_208_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9612" *) FpMul_8U_23U_lor_8_lpi_1_dfm_7;
  assign _05801_ = _05800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9612" *) _00978_;
  assign _05802_ = _00979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9613" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign _05803_ = _05413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9613" *) _00980_;
  assign _05804_ = _05791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9616" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign _05805_ = _05804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9616" *) _00766_;
  assign _05806_ = _05805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9616" *) FpMul_8U_23U_lor_8_lpi_1_dfm_6;
  assign _05807_ = _05806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9617" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _05808_ = _05807_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9617" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign _05809_ = _05808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9617" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05810_ = _05794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9619" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign _05811_ = _05810_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9619" *) _00766_;
  assign _05812_ = _05811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9620" *) FpMul_8U_23U_lor_8_lpi_1_dfm_6;
  assign _05813_ = _05812_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9620" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _05814_ = _05813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9620" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign _05815_ = _05814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9620" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05816_ = _05797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9625" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign _05817_ = _05816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9625" *) _00766_;
  assign _05818_ = _05817_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9626" *) FpMul_8U_23U_lor_8_lpi_1_dfm_6;
  assign _05819_ = _05818_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9626" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _05820_ = _05819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9626" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign _05821_ = _05820_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9626" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05822_ = nor_208_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9628" *) _00752_;
  assign _05823_ = _05822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9629" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _05824_ = _05823_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9629" *) mul_mul_land_3_lpi_1_dfm_6;
  assign _05825_ = _05824_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9629" *) IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  assign _05826_ = _05825_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9630" *) mul_mul_land_3_lpi_1_dfm_st_5;
  assign _05827_ = _05826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9630" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign _05828_ = _05827_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9630" *) FpMul_8U_23U_lor_8_lpi_1_dfm_7;
  assign _05829_ = _05828_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9630" *) _00978_;
  assign _05830_ = IsNaN_8U_23U_land_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9633" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign or_387_nl = _05830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9633" *) mul_mul_land_lpi_1_dfm_5;
  assign _05831_ = nor_190_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9634" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign _05832_ = _05831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9635" *) _00780_;
  assign _05833_ = _05832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9635" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign or_390_nl = _05833_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9635" *) mul_mul_land_lpi_1_dfm_5;
  assign _05834_ = _00981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9637" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign _05835_ = _05834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9638" *) _00780_;
  assign _05836_ = _05835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9638" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign or_391_nl = _05836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9638" *) mul_mul_land_lpi_1_dfm_5;
  assign _05837_ = _00982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9641" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign _05838_ = _05837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9642" *) _00780_;
  assign _05839_ = _05838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9642" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign or_395_nl = _05839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9642" *) mul_mul_land_lpi_1_dfm_5;
  assign _05840_ = _00634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9645" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm;
  assign or_828_nl = _00983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9646" *) mux_131_nl;
  assign _05841_ = or_435_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9650" *) mux_133_nl;
  assign or_424_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9651" *) _00984_;
  assign _05842_ = nor_193_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9656" *) mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2;
  assign _05843_ = _05436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9661" *) mux_135_nl;
  assign _05844_ = _00779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9664" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05845_ = _05844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9664" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05846_ = _05845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9664" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign _05847_ = _05846_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9664" *) not_tmp_121;
  assign _05848_ = _00986_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9666" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05849_ = _05848_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9666" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05850_ = _05849_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9667" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign _05851_ = _05850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9667" *) not_tmp_121;
  assign _05852_ = or_tmp_173 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9670" *) mul_mul_land_lpi_1_dfm_st_5;
  assign _05853_ = _05852_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9670" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_4;
  assign _05854_ = _05853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9671" *) _00987_;
  assign _05855_ = nor_190_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9673" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _05856_ = _05855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9674" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign or_414_nl = _05856_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9674" *) mul_mul_land_lpi_1_dfm_5;
  assign _05857_ = _00981_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9676" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _05858_ = _05857_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9676" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign or_415_nl = _05858_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9676" *) mul_mul_land_lpi_1_dfm_5;
  assign _05859_ = _00982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9679" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _05860_ = _05859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9680" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign or_418_nl = _05860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9680" *) mul_mul_land_lpi_1_dfm_5;
  assign _05861_ = _05339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9685" *) mux_142_nl;
  assign _05862_ = _00988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9687" *) _00752_;
  assign _05863_ = _05862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9687" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _05864_ = _05863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9688" *) mul_mul_land_lpi_1_dfm_6;
  assign _05865_ = _05864_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9688" *) IsNaN_8U_23U_land_lpi_1_dfm_8;
  assign _05866_ = _05865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9688" *) mul_mul_land_lpi_1_dfm_st_5;
  assign _05867_ = _05866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9689" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _05868_ = _05867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9689" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_4;
  assign _05869_ = _05868_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9689" *) _00984_;
  assign or_429_nl = or_430_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9692" *) or_tmp_411;
  assign or_436_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9697" *) or_tmp_411;
  assign _05870_ = io_read_cfg_mul_bypass_rsc_svs_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9701" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign _05871_ = _05870_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9701" *) mul_mul_land_lpi_1_dfm_5;
  assign _05872_ = nor_170_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9702" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05873_ = _05872_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9703" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign _05874_ = _05873_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9703" *) mul_mul_land_lpi_1_dfm_5;
  assign _05875_ = FpMul_8U_23U_p_mant_p1_sva[47] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9705" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05876_ = _05875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9705" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign _05877_ = _05876_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9705" *) mul_mul_land_lpi_1_dfm_5;
  assign _05878_ = _00989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9710" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05879_ = _05878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9710" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign or_453_nl = _05879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9710" *) mul_mul_land_lpi_1_dfm_5;
  assign _05880_ = FpMul_8U_23U_lor_1_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9712" *) mux_154_nl;
  assign _05881_ = nor_174_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9718" *) FpMul_8U_23U_lor_1_lpi_1_dfm_7;
  assign _05882_ = _05881_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9718" *) _00991_;
  assign _05883_ = _00992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9719" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _05884_ = _05436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9719" *) _00993_;
  assign _05885_ = _05872_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9722" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05886_ = _05885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9722" *) _00766_;
  assign _05887_ = _05886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9722" *) FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  assign _05888_ = _05887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9723" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _05889_ = _05888_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9723" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign _05890_ = _05889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9723" *) mul_mul_land_lpi_1_dfm_5;
  assign _05891_ = _05875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9725" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05892_ = _05891_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9725" *) _00766_;
  assign _05893_ = _05892_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9726" *) FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  assign _05894_ = _05893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9726" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _05895_ = _05894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9726" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign _05896_ = _05895_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9726" *) mul_mul_land_lpi_1_dfm_5;
  assign _05897_ = _05878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9731" *) mul_mul_land_lpi_1_dfm_st_4;
  assign _05898_ = _05897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9731" *) _00766_;
  assign _05899_ = _05898_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9732" *) FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  assign _05900_ = _05899_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9732" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _05901_ = _05900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9732" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign _05902_ = _05901_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9732" *) mul_mul_land_lpi_1_dfm_5;
  assign _05903_ = nor_174_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9734" *) _00752_;
  assign _05904_ = _05903_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9735" *) io_read_cfg_mul_bypass_rsc_svs_5;
  assign _05905_ = _05904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9735" *) mul_mul_land_lpi_1_dfm_6;
  assign _05906_ = _05905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9735" *) IsNaN_8U_23U_land_lpi_1_dfm_8;
  assign _05907_ = _05906_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9736" *) mul_mul_land_lpi_1_dfm_st_5;
  assign _05908_ = _05907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9736" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _05909_ = _05908_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9736" *) FpMul_8U_23U_lor_1_lpi_1_dfm_7;
  assign _05910_ = _05909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9736" *) _00991_;
  assign _05911_ = mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9739" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign or_511_nl = _05911_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9739" *) or_tmp_167;
  assign _05912_ = _00767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9741" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign _05913_ = _05912_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9741" *) or_tmp_167;
  assign _05914_ = or_27_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9744" *) _00768_;
  assign or_509_nl = _05914_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9744" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  assign _05915_ = nor_143_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9752" *) or_27_cse;
  assign _05916_ = _05915_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9753" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05917_ = _05916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9753" *) mul_mul_land_1_lpi_1_dfm_st_4;
  assign _05918_ = _05917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9753" *) _00766_;
  assign _05919_ = or_744_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9758" *) mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign _05920_ = _05919_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9758" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign or_519_nl = _05920_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9758" *) or_tmp_167;
  assign _05921_ = or_744_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9761" *) _00771_;
  assign _05922_ = _05921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9761" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign _05923_ = _05922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9761" *) or_tmp_167;
  assign _05924_ = _05916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9771" *) mul_mul_land_2_lpi_1_dfm_st_4;
  assign _05925_ = _05924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9771" *) _00766_;
  assign _05926_ = or_745_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9776" *) mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign _05927_ = _05926_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9776" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign or_527_nl = _05927_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9776" *) or_tmp_167;
  assign _05928_ = or_745_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9779" *) _00775_;
  assign _05929_ = _05928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9779" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign _05930_ = _05929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9779" *) or_tmp_167;
  assign _05931_ = _05916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9789" *) mul_mul_land_3_lpi_1_dfm_st_4;
  assign _05932_ = _05931_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9789" *) _00766_;
  assign _05933_ = or_430_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9794" *) mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign or_535_nl = _05933_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9794" *) or_tmp_411;
  assign _05934_ = or_430_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9797" *) _00779_;
  assign _05935_ = _05934_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9797" *) or_tmp_411;
  assign _05936_ = FpMul_8U_23U_p_mant_p1_sva[47] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9801" *) _00994_;
  assign _05937_ = or_tmp_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9812" *) IsNaN_8U_23U_land_1_lpi_1_dfm_4;
  assign _05938_ = _05937_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9812" *) mul_mul_land_1_lpi_1_dfm_2;
  assign _05939_ = _00640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9814" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05940_ = _05939_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9814" *) mul_mul_land_1_lpi_1_dfm_st_1;
  assign _05941_ = _05940_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9815" *) IsNaN_8U_23U_land_1_lpi_1_dfm_4;
  assign _05942_ = _05941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9815" *) mul_mul_land_1_lpi_1_dfm_2;
  assign or_540_nl = or_27_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9816" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st_1;
  assign _05943_ = _05362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9819" *) _00765_;
  assign _05944_ = _05943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9820" *) chn_mul_out_rsci_bawt;
  assign _05945_ = _05944_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9820" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _05946_ = _05945_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9820" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign _05947_ = _05946_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9820" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05948_ = mul_mul_land_1_lpi_1_dfm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9823" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05949_ = or_74_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9825" *) mul_mul_land_1_lpi_1_dfm_5;
  assign _05950_ = _05949_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9825" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05951_ = _05950_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9825" *) _00766_;
  assign _05952_ = or_tmp_15 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9830" *) IsNaN_8U_23U_land_2_lpi_1_dfm_4;
  assign _05953_ = _05952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9830" *) mul_mul_land_2_lpi_1_dfm_2;
  assign _05954_ = _00641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9832" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05955_ = _05954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9832" *) mul_mul_land_2_lpi_1_dfm_st_1;
  assign _05956_ = _05955_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9833" *) IsNaN_8U_23U_land_2_lpi_1_dfm_4;
  assign _05957_ = _05956_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9833" *) mul_mul_land_2_lpi_1_dfm_2;
  assign or_551_nl = or_27_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9834" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st_1;
  assign _05958_ = _05385_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9837" *) _00765_;
  assign _05959_ = _05958_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9838" *) chn_mul_out_rsci_bawt;
  assign _05960_ = _05959_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9838" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _05961_ = _05960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9838" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign _05962_ = _05961_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9838" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05963_ = mul_mul_land_2_lpi_1_dfm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9841" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05964_ = or_74_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9843" *) mul_mul_land_2_lpi_1_dfm_5;
  assign _05965_ = _05964_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9843" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05966_ = _05965_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9843" *) _00766_;
  assign _05967_ = or_tmp_29 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9848" *) IsNaN_8U_23U_land_3_lpi_1_dfm_4;
  assign _05968_ = _05967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9848" *) mul_mul_land_3_lpi_1_dfm_2;
  assign _05969_ = _00642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9850" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05970_ = _05969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9850" *) mul_mul_land_3_lpi_1_dfm_st_1;
  assign _05971_ = _05970_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9851" *) IsNaN_8U_23U_land_3_lpi_1_dfm_4;
  assign _05972_ = _05971_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9851" *) mul_mul_land_3_lpi_1_dfm_2;
  assign or_561_nl = or_27_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9852" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st_1;
  assign _05973_ = _05408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9855" *) _00765_;
  assign _05974_ = _05973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9856" *) chn_mul_out_rsci_bawt;
  assign _05975_ = _05974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9856" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _05976_ = _05975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9856" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign _05977_ = _05976_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9856" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05978_ = mul_mul_land_3_lpi_1_dfm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9859" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05979_ = or_74_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9861" *) mul_mul_land_3_lpi_1_dfm_5;
  assign _05980_ = _05979_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9861" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05981_ = _05980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9861" *) _00766_;
  assign _05982_ = or_tmp_46 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9866" *) IsNaN_8U_23U_land_lpi_1_dfm_4;
  assign _05983_ = _05982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9866" *) mul_mul_land_lpi_1_dfm_2;
  assign _05984_ = _00643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9868" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05985_ = _05984_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9868" *) mul_mul_land_lpi_1_dfm_st_1;
  assign _05986_ = _05985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9869" *) IsNaN_8U_23U_land_lpi_1_dfm_4;
  assign _05987_ = _05986_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9869" *) mul_mul_land_lpi_1_dfm_2;
  assign or_571_nl = or_27_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9870" *) IsNaN_8U_23U_land_lpi_1_dfm_st_1;
  assign _05988_ = or_435_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9873" *) _00765_;
  assign _05989_ = _05988_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9874" *) chn_mul_out_rsci_bawt;
  assign _05990_ = _05989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9874" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _05991_ = _05990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9874" *) IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign _05992_ = _05991_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9874" *) mul_mul_land_lpi_1_dfm_5;
  assign _05993_ = mul_mul_land_lpi_1_dfm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9877" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _05994_ = or_74_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9879" *) mul_mul_land_lpi_1_dfm_5;
  assign _05995_ = _05994_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9879" *) io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _05996_ = _05995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9879" *) _00766_;
  assign _05997_ = or_tmp_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9881" *) nor_118_cse;
  assign or_473_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_st | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9883" *) _00995_;
  assign _05998_ = _00862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9886" *) mul_mul_land_1_lpi_1_dfm_st_1;
  assign _05999_ = _05998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9886" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _06000_ = _05999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9886" *) IsZero_8U_23U_land_1_lpi_1_dfm_4;
  assign _06001_ = _06000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9887" *) mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign or_474_nl = _06001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9887" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp;
  assign _06002_ = or_tmp_15 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9890" *) nor_117_cse;
  assign or_486_nl = FpMul_8U_23U_lor_7_lpi_1_dfm_st | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9892" *) _00996_;
  assign _06003_ = _00863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9895" *) mul_mul_land_2_lpi_1_dfm_st_1;
  assign _06004_ = _06003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9895" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _06005_ = _06004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9895" *) IsZero_8U_23U_land_2_lpi_1_dfm_4;
  assign _06006_ = _06005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9896" *) mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign or_487_nl = _06006_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9896" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp;
  assign _06007_ = or_tmp_29 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9899" *) nor_116_cse;
  assign or_494_nl = FpMul_8U_23U_lor_8_lpi_1_dfm_st | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9901" *) _00997_;
  assign _06008_ = _00864_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9904" *) mul_mul_land_3_lpi_1_dfm_st_1;
  assign _06009_ = _06008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9904" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _06010_ = _06009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9904" *) IsZero_8U_23U_land_3_lpi_1_dfm_4;
  assign _06011_ = _06010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9905" *) mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign or_495_nl = _06011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9905" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp;
  assign _06012_ = or_tmp_46 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9910" *) nor_115_cse;
  assign or_502_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9912" *) _00998_;
  assign _06013_ = _00865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9915" *) mul_mul_land_lpi_1_dfm_st_1;
  assign _06014_ = _06013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9915" *) io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _06015_ = _06014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9916" *) mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign _06016_ = _06015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9916" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp;
  assign or_503_nl = _06016_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9916" *) IsZero_8U_23U_land_lpi_1_dfm_4;
  assign _06017_ = _00644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *) _00648_;
  assign _06018_ = _00645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *) _00649_;
  assign _06019_ = _00646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *) _00650_;
  assign _06020_ = _00647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9936" *) _00651_;
  assign _06021_ = _06017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *) _00652_;
  assign _06022_ = _06018_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *) _00653_;
  assign _06023_ = _06019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *) _00654_;
  assign _06024_ = _06020_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9937" *) _00655_;
  assign _06025_ = _00656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *) _00660_;
  assign _06026_ = _00657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *) _00661_;
  assign _06027_ = _00658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *) _00662_;
  assign _06028_ = _00659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9949" *) _00663_;
  assign _06029_ = _06025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *) _00664_;
  assign _06030_ = _06026_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *) _00665_;
  assign _06031_ = _06027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *) _00666_;
  assign _06032_ = _06028_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9950" *) _00667_;
  assign _06033_ = _00668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *) _00672_;
  assign _06034_ = _00669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *) _00673_;
  assign _06035_ = _00670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *) _00674_;
  assign _06036_ = _00671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9962" *) _00675_;
  assign FpMul_8U_23U_o_mant_1_lpi_1_dfm_3 = _06033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *) _00676_;
  assign FpMul_8U_23U_o_mant_2_lpi_1_dfm_3 = _06034_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *) _00677_;
  assign FpMul_8U_23U_o_mant_3_lpi_1_dfm_3 = _06035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *) _00678_;
  assign FpMul_8U_23U_o_mant_lpi_1_dfm_3 = _06036_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9963" *) _00679_;
  assign _06037_ = _00680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *) _00684_;
  assign _06038_ = _00681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *) _00685_;
  assign _06039_ = _00682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *) _00686_;
  assign _06040_ = _00683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9976" *) _00687_;
  assign _06041_ = _06037_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *) _00688_;
  assign _06042_ = _06038_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *) _00689_;
  assign _06043_ = _06039_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *) _00690_;
  assign _06044_ = _06040_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9977" *) _00691_;
  assign _06045_ = _06041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *) _00692_;
  assign _06046_ = _06042_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *) _00693_;
  assign _06047_ = _06043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *) _00694_;
  assign _06048_ = _06044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9978" *) _00695_;
  assign _06049_ = _00696_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *) _00700_;
  assign _06050_ = _00697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *) _00701_;
  assign _06051_ = _00698_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *) _00702_;
  assign _06052_ = _00699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9990" *) _00703_;
  assign FpMul_8U_23U_o_expo_1_lpi_1_dfm = _06049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *) _00704_;
  assign FpMul_8U_23U_o_expo_2_lpi_1_dfm = _06050_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *) _00705_;
  assign FpMul_8U_23U_o_expo_3_lpi_1_dfm = _06051_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *) _00706_;
  assign FpMul_8U_23U_o_expo_lpi_1_dfm = _06052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9991" *) _00707_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm <= _00277_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= 1'b0;
    else
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= _00273_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm <= _00261_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= 1'b0;
    else
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= _00257_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm <= _00245_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= 1'b0;
    else
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= _00241_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm <= _00229_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= 1'b0;
    else
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs <= _00225_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_mul_src_1_sva_st <= 1'b0;
    else
      cfg_mul_src_1_sva_st <= _00172_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_lpi_1_dfm <= 1'b0;
    else
      IsZero_8U_23U_land_lpi_1_dfm <= _00164_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_st <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_st <= _00143_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_3_lpi_1_dfm <= 1'b0;
    else
      IsZero_8U_23U_land_3_lpi_1_dfm <= _00161_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_st <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_st <= _00136_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_2_lpi_1_dfm <= 1'b0;
    else
      IsZero_8U_23U_land_2_lpi_1_dfm <= _00158_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_st <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_st <= _00129_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_1_lpi_1_dfm <= 1'b0;
    else
      IsZero_8U_23U_land_1_lpi_1_dfm <= _00155_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_st <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_st <= _00122_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_1_lpi_1_dfm_st <= 1'b0;
    else
      FpMul_8U_23U_lor_1_lpi_1_dfm_st <= _00065_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_1_land_lpi_1_dfm_5 <= 1'b0;
    else
      IsZero_8U_23U_1_land_lpi_1_dfm_5 <= _00153_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_8_lpi_1_dfm_st <= 1'b0;
    else
      FpMul_8U_23U_lor_8_lpi_1_dfm_st <= _00080_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_1_land_3_lpi_1_dfm_5 <= 1'b0;
    else
      IsZero_8U_23U_1_land_3_lpi_1_dfm_5 <= _00151_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_7_lpi_1_dfm_st <= 1'b0;
    else
      FpMul_8U_23U_lor_7_lpi_1_dfm_st <= _00075_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_1_land_2_lpi_1_dfm_5 <= 1'b0;
    else
      IsZero_8U_23U_1_land_2_lpi_1_dfm_5 <= _00149_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_6_lpi_1_dfm_st <= 1'b0;
    else
      FpMul_8U_23U_lor_6_lpi_1_dfm_st <= _00070_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_1_land_1_lpi_1_dfm_5 <= 1'b0;
    else
      IsZero_8U_23U_1_land_1_lpi_1_dfm_5 <= _00147_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <= 1'b0;
    else
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <= _00274_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_mant_p1_sva <= 48'b000000000000000000000000000000000000000000000000;
    else
      FpMul_8U_23U_p_mant_p1_sva <= _00102_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <= 1'b0;
    else
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <= _00258_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_mant_p1_3_sva <= 48'b000000000000000000000000000000000000000000000000;
    else
      FpMul_8U_23U_p_mant_p1_3_sva <= _00101_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <= 1'b0;
    else
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <= _00242_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_mant_p1_2_sva <= 48'b000000000000000000000000000000000000000000000000;
    else
      FpMul_8U_23U_p_mant_p1_2_sva <= _00100_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_truncate_1_sva_3 <= 10'b0000000000;
    else
      cfg_truncate_1_sva_3 <= _00175_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <= 1'b0;
    else
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 <= _00226_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_mant_p1_1_sva <= 48'b000000000000000000000000000000000000000000000000;
    else
      FpMul_8U_23U_p_mant_p1_1_sva <= _00099_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_mux_49_itm_3 <= 1'b0;
    else
      FpMul_8U_23U_mux_49_itm_3 <= _00089_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_lpi_1_dfm_6 <= _00117_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_1_lpi_1_dfm_6 <= 1'b0;
    else
      FpMul_8U_23U_lor_1_lpi_1_dfm_6 <= _00063_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_mux_36_itm_3 <= 1'b0;
    else
      FpMul_8U_23U_mux_36_itm_3 <= _00087_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 <= _00115_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_8_lpi_1_dfm_6 <= 1'b0;
    else
      FpMul_8U_23U_lor_8_lpi_1_dfm_6 <= _00078_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_mux_23_itm_3 <= 1'b0;
    else
      FpMul_8U_23U_mux_23_itm_3 <= _00085_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 <= _00113_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_7_lpi_1_dfm_6 <= 1'b0;
    else
      FpMul_8U_23U_lor_7_lpi_1_dfm_6 <= _00073_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_mux_10_itm_3 <= 1'b0;
    else
      FpMul_8U_23U_mux_10_itm_3 <= _00083_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 <= _00111_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_6_lpi_1_dfm_6 <= 1'b0;
    else
      FpMul_8U_23U_lor_6_lpi_1_dfm_6 <= _00068_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= 1'b0;
    else
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= _00281_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= 1'b0;
    else
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= _00279_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_48U_24U_else_carry_sva <= 1'b0;
    else
      FpMantRNE_48U_24U_else_carry_sva <= _00037_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_FpMul_8U_23U_and_14_itm <= 1'b0;
    else
      FpMul_8U_23U_FpMul_8U_23U_and_14_itm <= _00043_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st <= 1'b0;
    else
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st <= _00268_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm <= 23'b00000000000000000000000;
    else
      else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm <= _00210_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_3_30_23_5_itm <= 8'b00000000;
    else
      else_MulOp_data_slc_else_MulOp_data_3_30_23_5_itm <= _00212_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_expo_sva_1 <= 8'b00000000;
    else
      FpMul_8U_23U_p_expo_sva_1 <= _00097_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm <= _00051_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= 1'b0;
    else
      mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= _00271_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 <= 23'b00000000000000000000000;
    else
      mul_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 <= _00270_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2 <= _00061_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= 1'b0;
    else
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= _00265_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= 1'b0;
    else
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= _00263_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_48U_24U_else_carry_3_sva <= 1'b0;
    else
      FpMantRNE_48U_24U_else_carry_3_sva <= _00035_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_FpMul_8U_23U_and_13_itm <= 1'b0;
    else
      FpMul_8U_23U_FpMul_8U_23U_and_13_itm <= _00041_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st <= 1'b0;
    else
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st <= _00252_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm <= 23'b00000000000000000000000;
    else
      else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm <= _00207_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_2_30_23_5_itm <= 8'b00000000;
    else
      else_MulOp_data_slc_else_MulOp_data_2_30_23_5_itm <= _00209_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_expo_3_sva_1 <= 8'b00000000;
    else
      FpMul_8U_23U_p_expo_3_sva_1 <= _00095_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm <= _00049_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= 1'b0;
    else
      mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= _00255_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 <= 23'b00000000000000000000000;
    else
      mul_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 <= _00254_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2 <= _00059_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= 1'b0;
    else
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= _00249_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= 1'b0;
    else
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= _00247_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_48U_24U_else_carry_2_sva <= 1'b0;
    else
      FpMantRNE_48U_24U_else_carry_2_sva <= _00033_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_FpMul_8U_23U_and_12_itm <= 1'b0;
    else
      FpMul_8U_23U_FpMul_8U_23U_and_12_itm <= _00039_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st <= 1'b0;
    else
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st <= _00236_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm <= 23'b00000000000000000000000;
    else
      else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm <= _00204_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_1_30_23_5_itm <= 8'b00000000;
    else
      else_MulOp_data_slc_else_MulOp_data_1_30_23_5_itm <= _00206_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_expo_2_sva_1 <= 8'b00000000;
    else
      FpMul_8U_23U_p_expo_2_sva_1 <= _00093_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm <= _00047_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= 1'b0;
    else
      mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= _00239_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 <= 23'b00000000000000000000000;
    else
      mul_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 <= _00238_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2 <= _00057_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= 1'b0;
    else
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm <= _00233_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= 1'b0;
    else
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm <= _00231_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_48U_24U_else_carry_1_sva <= 1'b0;
    else
      FpMantRNE_48U_24U_else_carry_1_sva <= _00031_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_FpMul_8U_23U_and_itm <= 1'b0;
    else
      FpMul_8U_23U_FpMul_8U_23U_and_itm <= _00045_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st <= 1'b0;
    else
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st <= _00220_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm <= 23'b00000000000000000000000;
    else
      else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm <= _00201_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_0_30_23_5_itm <= 8'b00000000;
    else
      else_MulOp_data_slc_else_MulOp_data_0_30_23_5_itm <= _00203_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_expo_1_sva_1 <= 8'b00000000;
    else
      FpMul_8U_23U_p_expo_1_sva_1 <= _00091_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm <= _00053_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= 1'b0;
    else
      mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm <= _00223_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 <= 23'b00000000000000000000000;
    else
      mul_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1 <= _00222_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2 <= _00055_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_mul_src_1_sva_st_1 <= 1'b0;
    else
      cfg_mul_src_1_sva_st_1 <= _00173_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_1_lpi_1_dfm_st_1 <= 1'b0;
    else
      mul_mul_land_1_lpi_1_dfm_st_1 <= _00286_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_2_lpi_1_dfm_st_1 <= 1'b0;
    else
      mul_mul_land_2_lpi_1_dfm_st_1 <= _00292_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_3_lpi_1_dfm_st_1 <= 1'b0;
    else
      mul_mul_land_3_lpi_1_dfm_st_1 <= _00298_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_lpi_1_dfm_st_1 <= 1'b0;
    else
      mul_mul_land_lpi_1_dfm_st_1 <= _00304_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_lpi_1_dfm_4 <= 1'b0;
    else
      IsZero_8U_23U_land_lpi_1_dfm_4 <= _00165_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_st_1 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_st_1 <= _00144_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_3_lpi_1_dfm_4 <= 1'b0;
    else
      IsZero_8U_23U_land_3_lpi_1_dfm_4 <= _00162_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_1 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_1 <= _00137_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_2_lpi_1_dfm_4 <= 1'b0;
    else
      IsZero_8U_23U_land_2_lpi_1_dfm_4 <= _00159_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_1 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_1 <= _00130_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_mul_src_1_sva_1 <= 1'b0;
    else
      cfg_mul_src_1_sva_1 <= _00171_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_mul_op_1_sva_1 <= 32'd0;
    else
      cfg_mul_op_1_sva_1 <= _00170_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_1_lpi_1_dfm_4 <= 1'b0;
    else
      IsZero_8U_23U_land_1_lpi_1_dfm_4 <= _00156_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_1 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_1 <= _00123_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_4 <= _00140_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_4 <= _00133_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_4 <= _00126_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_4 <= _00119_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      io_read_cfg_mul_bypass_rsc_svs_st_1 <= 1'b0;
    else
      io_read_cfg_mul_bypass_rsc_svs_st_1 <= _00214_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_1_lpi_1_dfm_2 <= 1'b0;
    else
      mul_mul_land_1_lpi_1_dfm_2 <= _00283_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_2_lpi_1_dfm_2 <= 1'b0;
    else
      mul_mul_land_2_lpi_1_dfm_2 <= _00289_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_3_lpi_1_dfm_2 <= 1'b0;
    else
      mul_mul_land_3_lpi_1_dfm_2 <= _00295_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_lpi_1_dfm_2 <= 1'b0;
    else
      mul_mul_land_lpi_1_dfm_2 <= _00301_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_truncate_1_sva_1 <= 10'b0000000000;
    else
      cfg_truncate_1_sva_1 <= _00174_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      MulIn_data_sva_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      MulIn_data_sva_1 <= _00169_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_1 <= 1'b0;
    else
      main_stage_v_1 <= _00216_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_1_lpi_1_dfm_st_5 <= 1'b0;
    else
      mul_mul_land_1_lpi_1_dfm_st_5 <= _00288_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_2_lpi_1_dfm_st_5 <= 1'b0;
    else
      mul_mul_land_2_lpi_1_dfm_st_5 <= _00294_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_3_lpi_1_dfm_st_5 <= 1'b0;
    else
      mul_mul_land_3_lpi_1_dfm_st_5 <= _00300_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_lpi_1_dfm_st_5 <= 1'b0;
    else
      mul_mul_land_lpi_1_dfm_st_5 <= _00306_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= 1'b0;
    else
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= _00282_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= 1'b0;
    else
      mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= _00280_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_48U_24U_else_carry_sva_2 <= 1'b0;
    else
      FpMantRNE_48U_24U_else_carry_sva_2 <= _00038_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    else
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2 <= _00269_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_1_lpi_1_dfm_7 <= 1'b0;
    else
      FpMul_8U_23U_lor_1_lpi_1_dfm_7 <= _00064_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 <= 1'b0;
    else
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 <= _00067_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_st_5 <= _00146_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm_2 <= 23'b00000000000000000000000;
    else
      else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm_2 <= _00211_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    else
      mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2 <= _00267_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2 <= 1'b0;
    else
      FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2 <= _00044_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= _00118_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_64_1 <= 1'b0;
    else
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_64_1 <= _00110_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 <= 1'b0;
    else
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 <= _00276_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= 1'b0;
    else
      mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= _00272_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2 <= _00052_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_3 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_3 <= _00062_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_expo_sva_5 <= 8'b00000000;
    else
      FpMul_8U_23U_p_expo_sva_5 <= _00098_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= 1'b0;
    else
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= _00266_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= 1'b0;
    else
      mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= _00264_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_48U_24U_else_carry_3_sva_2 <= 1'b0;
    else
      FpMantRNE_48U_24U_else_carry_3_sva_2 <= _00036_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    else
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2 <= _00253_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_8_lpi_1_dfm_7 <= 1'b0;
    else
      FpMul_8U_23U_lor_8_lpi_1_dfm_7 <= _00079_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 <= _00139_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_8_lpi_1_dfm_st_4 <= 1'b0;
    else
      FpMul_8U_23U_lor_8_lpi_1_dfm_st_4 <= _00082_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm_2 <= 23'b00000000000000000000000;
    else
      else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm_2 <= _00208_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    else
      mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2 <= _00251_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2 <= 1'b0;
    else
      FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2 <= _00042_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= _00116_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_64_1 <= 1'b0;
    else
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_64_1 <= _00108_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 <= 1'b0;
    else
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 <= _00260_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= 1'b0;
    else
      mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= _00256_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2 <= _00050_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_3 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_3 <= _00060_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_expo_3_sva_5 <= 8'b00000000;
    else
      FpMul_8U_23U_p_expo_3_sva_5 <= _00096_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= 1'b0;
    else
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= _00250_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= 1'b0;
    else
      mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= _00248_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_48U_24U_else_carry_2_sva_2 <= 1'b0;
    else
      FpMantRNE_48U_24U_else_carry_2_sva_2 <= _00034_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    else
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2 <= _00237_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_7_lpi_1_dfm_7 <= 1'b0;
    else
      FpMul_8U_23U_lor_7_lpi_1_dfm_7 <= _00074_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 <= _00132_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_7_lpi_1_dfm_st_4 <= 1'b0;
    else
      FpMul_8U_23U_lor_7_lpi_1_dfm_st_4 <= _00077_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm_2 <= 23'b00000000000000000000000;
    else
      else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm_2 <= _00205_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    else
      mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2 <= _00235_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2 <= 1'b0;
    else
      FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2 <= _00040_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= _00114_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_64_1 <= 1'b0;
    else
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_64_1 <= _00106_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 <= 1'b0;
    else
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 <= _00244_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= 1'b0;
    else
      mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= _00240_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2 <= _00048_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_3 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_3 <= _00058_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_expo_2_sva_5 <= 8'b00000000;
    else
      FpMul_8U_23U_p_expo_2_sva_5 <= _00094_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= 1'b0;
    else
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2 <= _00234_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= 1'b0;
    else
      mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2 <= _00232_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_48U_24U_else_carry_1_sva_2 <= 1'b0;
    else
      FpMantRNE_48U_24U_else_carry_1_sva_2 <= _00032_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2 <= 1'b0;
    else
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2 <= _00221_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_6_lpi_1_dfm_7 <= 1'b0;
    else
      FpMul_8U_23U_lor_6_lpi_1_dfm_7 <= _00069_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 <= _00125_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 <= 1'b0;
    else
      FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 <= _00072_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm_2 <= 23'b00000000000000000000000;
    else
      else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm_2 <= _00202_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_FpMul_8U_23U_and_itm_2 <= 1'b0;
    else
      FpMul_8U_23U_FpMul_8U_23U_and_itm_2 <= _00046_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2 <= 1'b0;
    else
      mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2 <= _00219_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= _00112_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_64_1 <= 1'b0;
    else
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_64_1 <= _00104_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 <= 1'b0;
    else
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4 <= _00228_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= 1'b0;
    else
      mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2 <= _00224_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2 <= _00054_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_3 <= 1'b0;
    else
      FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_3 <= _00056_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_p_expo_1_sva_5 <= 8'b00000000;
    else
      FpMul_8U_23U_p_expo_1_sva_5 <= _00092_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_mux_49_itm_4 <= 1'b0;
    else
      FpMul_8U_23U_mux_49_itm_4 <= _00090_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1 <= 32'd0;
    else
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1 <= _00109_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_mux_36_itm_4 <= 1'b0;
    else
      FpMul_8U_23U_mux_36_itm_4 <= _00088_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1 <= 32'd0;
    else
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1 <= _00107_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_mux_23_itm_4 <= 1'b0;
    else
      FpMul_8U_23U_mux_23_itm_4 <= _00086_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1 <= 32'd0;
    else
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1 <= _00105_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_mux_10_itm_4 <= 1'b0;
    else
      FpMul_8U_23U_mux_10_itm_4 <= _00084_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1 <= 32'd0;
    else
      IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1 <= _00103_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_8 <= _00142_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_8 <= _00135_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_8 <= _00128_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_8 <= _00121_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      io_read_cfg_mul_bypass_rsc_svs_5 <= 1'b0;
    else
      io_read_cfg_mul_bypass_rsc_svs_5 <= _00213_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_1_lpi_1_dfm_6 <= 1'b0;
    else
      mul_mul_land_1_lpi_1_dfm_6 <= _00285_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_2_lpi_1_dfm_6 <= 1'b0;
    else
      mul_mul_land_2_lpi_1_dfm_6 <= _00291_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_3_lpi_1_dfm_6 <= 1'b0;
    else
      mul_mul_land_3_lpi_1_dfm_6 <= _00297_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_lpi_1_dfm_6 <= 1'b0;
    else
      mul_mul_land_lpi_1_dfm_6 <= _00303_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      MulIn_data_sva_133 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      MulIn_data_sva_133 <= _00168_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_3 <= 1'b0;
    else
      main_stage_v_3 <= _00218_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_1_lpi_1_dfm_st_4 <= 1'b0;
    else
      mul_mul_land_1_lpi_1_dfm_st_4 <= _00287_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_2_lpi_1_dfm_st_4 <= 1'b0;
    else
      mul_mul_land_2_lpi_1_dfm_st_4 <= _00293_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_3_lpi_1_dfm_st_4 <= 1'b0;
    else
      mul_mul_land_3_lpi_1_dfm_st_4 <= _00299_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_lpi_1_dfm_st_4 <= 1'b0;
    else
      mul_mul_land_lpi_1_dfm_st_4 <= _00305_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 <= 1'b0;
    else
      FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 <= _00066_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_2 <= _00278_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 <= 1'b0;
    else
      mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 <= _00275_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_st_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_st_4 <= _00145_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_3_lpi_1_dfm_2_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      else_MulOp_data_3_lpi_1_dfm_2_30_0_1 <= _00200_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_1_land_lpi_1_dfm_6 <= 1'b0;
    else
      IsZero_8U_23U_1_land_lpi_1_dfm_6 <= _00154_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_lpi_1_dfm_6 <= 1'b0;
    else
      IsZero_8U_23U_land_lpi_1_dfm_6 <= _00166_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_2 <= _00262_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 <= 1'b0;
    else
      FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 <= _00081_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 <= 1'b0;
    else
      mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 <= _00259_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 <= _00138_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_2_lpi_1_dfm_2_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      else_MulOp_data_2_lpi_1_dfm_2_30_0_1 <= _00199_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_1_land_3_lpi_1_dfm_6 <= 1'b0;
    else
      IsZero_8U_23U_1_land_3_lpi_1_dfm_6 <= _00152_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_3_lpi_1_dfm_6 <= 1'b0;
    else
      IsZero_8U_23U_land_3_lpi_1_dfm_6 <= _00163_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_2 <= _00246_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 <= 1'b0;
    else
      FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 <= _00076_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 <= 1'b0;
    else
      mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 <= _00243_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 <= _00131_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_1_lpi_1_dfm_2_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      else_MulOp_data_1_lpi_1_dfm_2_30_0_1 <= _00198_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_1_land_2_lpi_1_dfm_6 <= 1'b0;
    else
      IsZero_8U_23U_1_land_2_lpi_1_dfm_6 <= _00150_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_2_lpi_1_dfm_6 <= 1'b0;
    else
      IsZero_8U_23U_land_2_lpi_1_dfm_6 <= _00160_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_2 <= _00230_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 <= 1'b0;
    else
      FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 <= _00071_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 <= 1'b0;
    else
      mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 <= _00227_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 <= _00124_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      else_MulOp_data_0_lpi_1_dfm_2_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      else_MulOp_data_0_lpi_1_dfm_2_30_0_1 <= _00197_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_1_land_1_lpi_1_dfm_6 <= 1'b0;
    else
      IsZero_8U_23U_1_land_1_lpi_1_dfm_6 <= _00148_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_1_lpi_1_dfm_5 <= 1'b0;
    else
      mul_mul_land_1_lpi_1_dfm_5 <= _00284_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_2_lpi_1_dfm_5 <= 1'b0;
    else
      mul_mul_land_2_lpi_1_dfm_5 <= _00290_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_3_lpi_1_dfm_5 <= 1'b0;
    else
      mul_mul_land_3_lpi_1_dfm_5 <= _00296_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mul_mul_land_lpi_1_dfm_5 <= 1'b0;
    else
      mul_mul_land_lpi_1_dfm_5 <= _00302_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_land_lpi_1_dfm_7 <= _00141_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_3_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_land_3_lpi_1_dfm_7 <= _00134_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_2_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_land_2_lpi_1_dfm_7 <= _00127_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_land_1_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_land_1_lpi_1_dfm_7 <= _00120_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      MulIn_data_sva_132 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      MulIn_data_sva_132 <= _00167_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      io_read_cfg_mul_bypass_rsc_svs_st_4 <= 1'b0;
    else
      io_read_cfg_mul_bypass_rsc_svs_st_4 <= _00215_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsZero_8U_23U_land_1_lpi_1_dfm_6 <= 1'b0;
    else
      IsZero_8U_23U_land_1_lpi_1_dfm_6 <= _00157_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_2 <= 1'b0;
    else
      main_stage_v_2 <= _00217_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_op_rsci_ld_core_psct <= 1'b0;
    else
      chn_mul_op_rsci_ld_core_psct <= _00179_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_chn_mul_out_rsci_ld_core_psct_cse <= 1'b0;
    else
      reg_chn_mul_out_rsci_ld_core_psct_cse <= _00308_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_126_119 <= 8'b00000000;
    else
      chn_mul_out_rsci_d_126_119 <= _00182_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_118_97 <= 22'b0000000000000000000000;
    else
      chn_mul_out_rsci_d_118_97 <= _00181_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_94_87 <= 8'b00000000;
    else
      chn_mul_out_rsci_d_94_87 <= _00193_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_86_65 <= 22'b0000000000000000000000;
    else
      chn_mul_out_rsci_d_86_65 <= _00192_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_62_55 <= 8'b00000000;
    else
      chn_mul_out_rsci_d_62_55 <= _00189_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_54_33 <= 22'b0000000000000000000000;
    else
      chn_mul_out_rsci_d_54_33 <= _00188_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_30_23 <= 8'b00000000;
    else
      chn_mul_out_rsci_d_30_23 <= _00185_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_22_1 <= 22'b0000000000000000000000;
    else
      chn_mul_out_rsci_d_22_1 <= _00184_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_127 <= 1'b0;
    else
      chn_mul_out_rsci_d_127 <= _00183_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_96 <= 1'b0;
    else
      chn_mul_out_rsci_d_96 <= _00195_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_95 <= 1'b0;
    else
      chn_mul_out_rsci_d_95 <= _00194_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_64 <= 1'b0;
    else
      chn_mul_out_rsci_d_64 <= _00191_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_63 <= 1'b0;
    else
      chn_mul_out_rsci_d_63 <= _00190_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_32 <= 1'b0;
    else
      chn_mul_out_rsci_d_32 <= _00187_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_31 <= 1'b0;
    else
      chn_mul_out_rsci_d_31 <= _00186_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_d_0 <= 1'b0;
    else
      chn_mul_out_rsci_d_0 <= _00180_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_in_rsci_ld_core_psct <= 1'b0;
    else
      chn_mul_in_rsci_ld_core_psct <= _00177_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_out_rsci_iswt0 <= 1'b0;
    else
      chn_mul_out_rsci_iswt0 <= _00196_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_op_rsci_iswt0 <= 1'b0;
    else
      chn_mul_op_rsci_iswt0 <= _00178_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_mul_in_rsci_iswt0 <= 1'b0;
    else
      chn_mul_in_rsci_iswt0 <= _00176_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
    else
      reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse <= _00307_;
  assign mux_182_nl = or_468_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_498_nl : mux_181_nl;
  assign mux_181_nl = mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_180_nl : or_503_nl;
  assign mux_180_nl = mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_179_nl : or_502_nl;
  assign mux_179_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_51 : nor_153_nl;
  assign mux_177_nl = or_468_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_490_cse : mux_176_nl;
  assign mux_176_nl = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_175_nl : or_495_nl;
  assign mux_175_nl = mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_174_nl : or_494_nl;
  assign mux_174_nl = FpMul_8U_23U_lor_8_lpi_1_dfm_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_40 : nor_155_nl;
  assign mux_172_nl = or_468_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_482_cse : mux_171_nl;
  assign mux_171_nl = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_170_nl : or_487_nl;
  assign mux_170_nl = mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_169_nl : or_486_nl;
  assign mux_169_nl = FpMul_8U_23U_lor_7_lpi_1_dfm_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_26 : nor_157_nl;
  assign mux_164_nl = or_468_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_469_cse : mux_163_nl;
  assign mux_163_nl = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_162_nl : or_474_nl;
  assign mux_162_nl = mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_161_nl : or_473_nl;
  assign mux_161_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_12 : nor_159_nl;
  assign mux_225_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_119_nl : nor_120_nl;
  assign mux_221_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_220_nl : nor_123_nl;
  assign mux_220_nl = or_571_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_121_nl : nor_122_nl;
  assign FpMul_8U_23U_oelse_1_mux_23_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_lor_1_lpi_1_dfm_mx0w0 : FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  assign mux_219_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_124_nl : nor_125_nl;
  assign mux_215_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_214_nl : nor_128_nl;
  assign mux_214_nl = or_561_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_126_nl : nor_127_nl;
  assign FpMul_8U_23U_oelse_1_mux_22_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0 : FpMul_8U_23U_lor_8_lpi_1_dfm_6;
  assign mux_213_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_129_nl : nor_130_nl;
  assign mux_209_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_208_nl : nor_133_nl;
  assign mux_208_nl = or_551_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_131_nl : nor_132_nl;
  assign FpMul_8U_23U_oelse_1_mux_21_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0 : FpMul_8U_23U_lor_7_lpi_1_dfm_6;
  assign mux_207_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_134_nl : nor_135_nl;
  assign mux_203_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_202_nl : nor_138_nl;
  assign mux_202_nl = or_540_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_136_nl : nor_137_nl;
  assign FpMul_8U_23U_oelse_1_mux_20_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0 : FpMul_8U_23U_lor_6_lpi_1_dfm_6;
  assign mux_201_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_FpMul_8U_23U_and_14_itm : mux_200_nl;
  assign mux_200_nl = or_430_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_198_nl : mux_199_nl;
  assign mux_199_nl = and_328_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_517 : and_tmp_5;
  assign mux_198_nl = _05936_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) and_tmp_5 : or_tmp_517;
  assign mux_197_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm : mux_196_nl;
  assign mux_196_nl = mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_535_nl : nor_342_nl;
  assign mux_195_nl = _05932_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_FpMul_8U_23U_and_13_itm : and_41_nl;
  assign mux_194_nl = or_745_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) _00002_ : or_531_nl;
  assign mux_193_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm : mux_192_nl;
  assign mux_192_nl = mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_527_nl : nor_140_nl;
  assign mux_191_nl = _05925_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_FpMul_8U_23U_and_12_itm : and_40_nl;
  assign mux_190_nl = or_744_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) _00001_ : or_523_nl;
  assign mux_189_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm : mux_188_nl;
  assign mux_188_nl = mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_519_nl : nor_142_nl;
  assign mux_187_nl = _05918_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_FpMul_8U_23U_and_itm : and_39_nl;
  assign mux_186_nl = or_743_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) _00000_ : or_515_nl;
  assign mux_185_nl = or_509_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm : mux_184_nl;
  assign mux_184_nl = mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_511_nl : nor_144_nl;
  assign mux_159_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_158_nl : nor_165_nl;
  assign mux_158_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_164_nl : and_331_nl;
  assign mux_157_nl = or_430_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_163_nl : nor_161_nl;
  assign mux_156_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) and_332_nl : nor_172_nl;
  assign mux_155_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_167_nl : nor_168_nl;
  assign mux_154_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_453_nl : nand_36_nl;
  assign mux_153_nl = or_430_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_171_nl : nor_169_nl;
  assign mux_149_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_436_nl : mux_148_nl;
  assign mux_148_nl = FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_415 : mux_tmp_140;
  assign mux_147_nl = or_424_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_429_nl : mux_146_nl;
  assign mux_146_nl = or_430_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_415 : mux_tmp_140;
  assign mux_143_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_181_nl : nor_183_nl;
  assign mux_142_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_141_nl : mux_140_nl;
  assign mux_141_nl = mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_395 : or_418_nl;
  assign mux_140_nl = mul_mul_4_FpMantRNE_48U_24U_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_395 : mux_139_nl;
  assign mux_139_nl = mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_414_nl : or_415_nl;
  assign mux_138_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_137_nl : nor_188_nl;
  assign mux_137_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_187_nl : nor_186_nl;
  assign mux_136_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_189_nl : nor_192_nl;
  assign mux_135_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsNaN_8U_23U_land_lpi_1_dfm_st_5 : nand_34_nl;
  assign mux_134_nl = FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_194_nl : and_334_nl;
  assign mux_133_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_387_nl : mux_132_nl;
  assign mux_132_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_828_nl : mux_130_nl;
  assign mux_131_nl = mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_371 : or_395_nl;
  assign mux_130_nl = mul_mul_4_FpMantRNE_48U_24U_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_371 : mux_129_nl;
  assign mux_129_nl = mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_390_nl : or_391_nl;
  assign mux_128_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_127_nl : nor_199_nl;
  assign mux_127_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_198_nl : and_335_nl;
  assign mux_126_nl = or_745_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_197_nl : nor_195_nl;
  assign mux_124_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) and_336_nl : nor_206_nl;
  assign mux_123_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_201_nl : nor_202_nl;
  assign mux_122_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_372_nl : nand_29_nl;
  assign mux_121_nl = or_745_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_205_nl : nor_203_nl;
  assign mux_116_nl = FpMul_8U_23U_lor_8_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_350_nl : mux_115_nl;
  assign mux_115_nl = or_tmp_332 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_336 : mux_tmp_109;
  assign mux_113_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_216_nl : nor_217_nl;
  assign mux_112_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_218_nl : nor_220_nl;
  assign mux_111_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_110_nl : mux_109_nl;
  assign mux_110_nl = mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_315 : or_338_nl;
  assign mux_109_nl = mul_mul_3_FpMantRNE_48U_24U_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_315 : mux_108_nl;
  assign mux_108_nl = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_334_nl : or_335_nl;
  assign mux_107_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_106_nl : nor_225_nl;
  assign mux_106_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_224_nl : nor_223_nl;
  assign mux_105_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_226_nl : nor_229_nl;
  assign mux_104_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st_5 : nand_27_nl;
  assign mux_103_nl = FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_231_nl : and_338_nl;
  assign mux_102_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_307_nl : mux_101_nl;
  assign mux_101_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_829_nl : mux_99_nl;
  assign mux_100_nl = mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_291 : or_315_nl;
  assign mux_99_nl = mul_mul_3_FpMantRNE_48U_24U_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_291 : mux_98_nl;
  assign mux_98_nl = mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_310_nl : or_311_nl;
  assign mux_97_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_96_nl : nor_236_nl;
  assign mux_96_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_235_nl : and_339_nl;
  assign mux_95_nl = or_744_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_234_nl : nor_232_nl;
  assign mux_93_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) and_340_nl : nor_243_nl;
  assign mux_92_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_238_nl : nor_239_nl;
  assign mux_91_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_292_nl : nand_22_nl;
  assign mux_90_nl = or_744_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_242_nl : nor_240_nl;
  assign mux_85_nl = FpMul_8U_23U_lor_7_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_270_nl : mux_84_nl;
  assign mux_84_nl = or_tmp_252 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_256 : mux_tmp_78;
  assign mux_82_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_253_nl : nor_254_nl;
  assign mux_81_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_255_nl : nor_257_nl;
  assign mux_80_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_79_nl : mux_78_nl;
  assign mux_79_nl = mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_235 : or_258_nl;
  assign mux_78_nl = mul_mul_2_FpMantRNE_48U_24U_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_235 : mux_77_nl;
  assign mux_77_nl = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_254_nl : or_255_nl;
  assign mux_76_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_75_nl : nor_262_nl;
  assign mux_75_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_261_nl : nor_260_nl;
  assign mux_74_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_263_nl : nor_266_nl;
  assign mux_73_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st_5 : nand_20_nl;
  assign mux_72_nl = FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_268_nl : and_342_nl;
  assign mux_71_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_227_nl : mux_70_nl;
  assign mux_70_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_830_nl : mux_68_nl;
  assign mux_69_nl = mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_211 : or_235_nl;
  assign mux_68_nl = mul_mul_2_FpMantRNE_48U_24U_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_211 : mux_67_nl;
  assign mux_67_nl = mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_230_nl : or_231_nl;
  assign mux_66_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_65_nl : nor_273_nl;
  assign mux_65_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_272_nl : and_343_nl;
  assign mux_64_nl = or_743_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_271_nl : nor_269_nl;
  assign mux_63_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_275_nl : nor_279_nl;
  assign mux_62_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_123 : or_211_nl;
  assign mux_61_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_210_nl : nand_15_nl;
  assign mux_60_nl = or_743_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_278_nl : nor_276_nl;
  assign mux_55_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_181_nl : mux_54_nl;
  assign mux_54_nl = FpMul_8U_23U_lor_6_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_185_nl : mux_tmp_48;
  assign mux_50_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_290_nl : nor_291_nl;
  assign mux_49_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_292_nl : nor_294_nl;
  assign mux_48_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_47_nl : mux_46_nl;
  assign mux_47_nl = mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_146 : or_169_nl;
  assign mux_46_nl = mul_mul_1_FpMantRNE_48U_24U_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_146 : mux_45_nl;
  assign mux_45_nl = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_165_nl : or_166_nl;
  assign mux_44_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_43_nl : nor_298_nl;
  assign mux_43_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_297_nl : nor_296_nl;
  assign mux_42_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) and_344_nl : nor_303_nl;
  assign mux_41_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st_5 : or_153_nl;
  assign mux_40_nl = mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_132 : nor_304_nl;
  assign mux_39_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_299_nl : nor_300_nl;
  assign mux_38_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_831_nl : mux_36_nl;
  assign mux_37_nl = mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_123 : or_147_nl;
  assign mux_36_nl = mul_mul_1_FpMantRNE_48U_24U_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_123 : mux_35_nl;
  assign mux_35_nl = mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_142_nl : or_143_nl;
  assign mux_24_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_23_nl : or_70_nl;
  assign mux_23_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_67_nl : or_tmp_51;
  assign mux_19_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_18_nl : or_59_nl;
  assign mux_18_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_56_nl : or_tmp_40;
  assign mux_14_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_13_nl : or_45_nl;
  assign mux_13_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_42_nl : or_tmp_26;
  assign mux_9_nl = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_8_nl : or_31_nl;
  assign mux_8_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_28_nl : or_tmp_12;
  assign _00030_ = IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) 8'b11111111 : mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  assign _00029_ = _01197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1[30:23] : 8'b11111111;
  assign FpMul_8U_23U_FpMul_8U_23U_and_18_nl = FpMul_8U_23U_lor_2_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) 8'b00000000 : FpMul_8U_23U_o_expo_lpi_1_dfm;
  assign _00010_ = IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10034|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10033" *) 22'b1111111111111111111111 : mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  assign _00009_ = _01197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10034|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10033" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1[22:1] : 22'b1111111111111111111111;
  assign _00028_ = IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) 8'b11111111 : mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  assign _00027_ = _01195_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1[30:23] : 8'b11111111;
  assign FpMul_8U_23U_FpMul_8U_23U_and_17_nl = FpMul_8U_23U_lor_11_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) 8'b00000000 : FpMul_8U_23U_o_expo_3_lpi_1_dfm;
  assign _00008_ = IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_3_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10034|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10033" *) 22'b1111111111111111111111 : mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  assign _00007_ = _01195_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10034|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10033" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1[22:1] : 22'b1111111111111111111111;
  assign _00026_ = IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) 8'b11111111 : mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  assign _00025_ = _01193_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1[30:23] : 8'b11111111;
  assign FpMul_8U_23U_FpMul_8U_23U_and_16_nl = FpMul_8U_23U_lor_10_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) 8'b00000000 : FpMul_8U_23U_o_expo_2_lpi_1_dfm;
  assign _00006_ = IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_2_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10034|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10033" *) 22'b1111111111111111111111 : mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  assign _00005_ = _01193_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10034|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10033" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1[22:1] : 22'b1111111111111111111111;
  assign _00024_ = IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) 8'b11111111 : mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_5_nl;
  assign _00023_ = _01191_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1[30:23] : 8'b11111111;
  assign FpMul_8U_23U_FpMul_8U_23U_and_15_nl = FpMul_8U_23U_lor_9_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) 8'b00000000 : FpMul_8U_23U_o_expo_1_lpi_1_dfm;
  assign _00004_ = IntShiftRight_64U_10U_32U_obits_fixed_and_unfl_1_sva ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10034|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10033" *) 22'b1111111111111111111111 : mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  assign _00003_ = _01191_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10034|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10033" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1[22:1] : 22'b1111111111111111111111;
  assign mul_mul_mux_115_nl = mul_mul_land_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) MulIn_data_sva_133[127] : mul_mul_else_mux_104_nl;
  assign mul_mul_else_mux_104_nl = and_dcpl_37 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_mux_49_itm_4 : mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  assign mul_mul_mux_114_nl = mul_mul_land_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) MulIn_data_sva_133[96] : mul_mul_else_mux_107_nl;
  assign mul_mul_else_mux_107_nl = and_dcpl_37 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_o_mant_lpi_1_dfm_3[0] : mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  assign mul_mul_mux_113_nl = mul_mul_land_3_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) MulIn_data_sva_133[95] : mul_mul_else_mux_77_nl;
  assign mul_mul_else_mux_77_nl = and_dcpl_37 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_mux_36_itm_4 : mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  assign mul_mul_mux_112_nl = mul_mul_land_3_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) MulIn_data_sva_133[64] : mul_mul_else_mux_80_nl;
  assign mul_mul_else_mux_80_nl = and_dcpl_37 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_o_mant_3_lpi_1_dfm_3[0] : mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  assign mul_mul_mux_111_nl = mul_mul_land_2_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) MulIn_data_sva_133[63] : mul_mul_else_mux_50_nl;
  assign mul_mul_else_mux_50_nl = and_dcpl_37 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_mux_23_itm_4 : mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  assign mul_mul_mux_110_nl = mul_mul_land_2_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) MulIn_data_sva_133[32] : mul_mul_else_mux_53_nl;
  assign mul_mul_else_mux_53_nl = and_dcpl_37 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_o_mant_2_lpi_1_dfm_3[0] : mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  assign mul_mul_mux_109_nl = mul_mul_land_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) MulIn_data_sva_133[31] : mul_mul_else_mux_23_nl;
  assign mul_mul_else_mux_23_nl = and_dcpl_37 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_mux_10_itm_4 : mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_2_nl;
  assign mul_mul_mux_108_nl = mul_mul_land_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) MulIn_data_sva_133[0] : mul_mul_else_mux_26_nl;
  assign mul_mul_else_mux_26_nl = and_dcpl_37 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_o_mant_1_lpi_1_dfm_3[0] : mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_nl;
  assign not_tmp_130 = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_175_nl : nor_176_nl;
  assign not_tmp_129 = mul_mul_land_lpi_1_dfm_st_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_177_nl : mux_150_nl;
  assign mux_150_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_179_nl : nor_180_nl;
  assign mux_tmp_140 = mul_mul_land_lpi_1_dfm_st_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_411 : mux_144_nl;
  assign mux_144_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_435_nl : or_tmp_173;
  assign mux_125_itm = mul_mul_land_3_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_336 : mux_tmp_109;
  assign not_tmp_107 = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_209_nl : nor_210_nl;
  assign not_tmp_106 = mul_mul_land_3_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_211_nl : mux_118_nl;
  assign mux_118_nl = mul_mul_land_3_lpi_1_dfm_st_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_212_nl : mux_117_nl;
  assign mux_117_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_214_nl : nor_215_nl;
  assign mux_tmp_109 = mul_mul_land_3_lpi_1_dfm_st_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_167 : mux_tmp_46;
  assign mux_94_itm = mul_mul_land_2_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_256 : mux_tmp_78;
  assign not_tmp_82 = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_246_nl : nor_247_nl;
  assign not_tmp_81 = mul_mul_land_2_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_248_nl : mux_87_nl;
  assign mux_87_nl = mul_mul_land_2_lpi_1_dfm_st_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_249_nl : mux_86_nl;
  assign mux_86_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_251_nl : nor_252_nl;
  assign mux_tmp_78 = mul_mul_land_2_lpi_1_dfm_st_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_167 : mux_tmp_46;
  assign not_tmp_55 = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_283_nl : nor_284_nl;
  assign not_tmp_54 = mul_mul_land_1_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_285_nl : mux_57_nl;
  assign mux_57_nl = or_193_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_286_nl : mux_56_nl;
  assign mux_56_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_288_nl : nor_289_nl;
  assign mux_tmp_48 = mul_mul_land_1_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_187_nl : mux_52_nl;
  assign mux_52_nl = mul_mul_land_1_lpi_1_dfm_st_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_167 : mux_tmp_46;
  assign mux_tmp_46 = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_189_cse : or_tmp_173;
  assign mux_22_itm = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_46 : or_65_nl;
  assign not_tmp_15 = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mux_20_nl : nor_323_nl;
  assign mux_20_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_322_nl : nor_321_nl;
  assign mux_17_itm = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_29 : or_54_nl;
  assign not_tmp_12 = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_324_nl : nor_325_nl;
  assign mux_15_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_490_cse : or_48_nl;
  assign mux_12_itm = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_15 : or_40_nl;
  assign not_tmp_8 = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_326_nl : nor_327_nl;
  assign mux_10_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_482_cse : or_34_nl;
  assign mux_7_itm = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_tmp_1 : or_26_nl;
  assign not_tmp_2 = and_18_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_nl : nor_331_nl;
  assign mux_5_nl = or_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_469_cse : or_19_nl;
  assign else_mux_tmp_30_23 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) chn_mul_op_rsci_d_mxwt[30:23] : cfg_mul_op_1_sva_1[30:23];
  assign else_mux_1_tmp_30_23 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) chn_mul_op_rsci_d_mxwt[62:55] : cfg_mul_op_1_sva_1[30:23];
  assign else_mux_2_tmp_30_23 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) chn_mul_op_rsci_d_mxwt[94:87] : cfg_mul_op_1_sva_1[30:23];
  assign else_mux_3_tmp_30_23 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) chn_mul_op_rsci_d_mxwt[126:119] : cfg_mul_op_1_sva_1[30:23];
  assign FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0 = mux_236_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10102|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10101" *) FpMul_8U_23U_p_mant_p1_sva_mx1[46:1] : FpMul_8U_23U_p_mant_p1_sva_mx1[45:0];
  assign mux_236_nl = or_430_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_p_mant_p1_sva[47] : mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0 = mux_235_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10102|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10101" *) FpMul_8U_23U_p_mant_p1_3_sva_mx1[46:1] : FpMul_8U_23U_p_mant_p1_3_sva_mx1[45:0];
  assign mux_235_nl = or_745_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_p_mant_p1_3_sva[47] : mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0 = mux_234_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10102|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10101" *) FpMul_8U_23U_p_mant_p1_2_sva_mx1[46:1] : FpMul_8U_23U_p_mant_p1_2_sva_mx1[45:0];
  assign mux_234_nl = or_744_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_p_mant_p1_2_sva[47] : mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0 = mux_233_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10102|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10101" *) FpMul_8U_23U_p_mant_p1_1_sva_mx1[46:1] : FpMul_8U_23U_p_mant_p1_1_sva_mx1[45:0];
  assign mux_233_nl = or_743_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_p_mant_p1_1_sva[47] : mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign else_MulOp_data_3_lpi_1_dfm_mx1 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10085|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10084" *) chn_mul_op_rsci_d_mxwt[127:96] : cfg_mul_op_1_sva_1;
  assign else_MulOp_data_3_lpi_1_dfm_mx0_30_0 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10068|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10067" *) chn_mul_op_rsci_d_mxwt[126:96] : cfg_mul_op_1_sva_1[30:0];
  assign else_MulOp_data_2_lpi_1_dfm_mx1 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10085|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10084" *) chn_mul_op_rsci_d_mxwt[95:64] : cfg_mul_op_1_sva_1;
  assign else_MulOp_data_2_lpi_1_dfm_mx0_30_0 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10068|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10067" *) chn_mul_op_rsci_d_mxwt[94:64] : cfg_mul_op_1_sva_1[30:0];
  assign else_MulOp_data_1_lpi_1_dfm_mx1 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10085|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10084" *) chn_mul_op_rsci_d_mxwt[63:32] : cfg_mul_op_1_sva_1;
  assign else_MulOp_data_1_lpi_1_dfm_mx0_30_0 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10068|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10067" *) chn_mul_op_rsci_d_mxwt[62:32] : cfg_mul_op_1_sva_1[30:0];
  assign else_MulOp_data_0_lpi_1_dfm_mx1 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10085|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10084" *) chn_mul_op_rsci_d_mxwt[31:0] : cfg_mul_op_1_sva_1;
  assign else_MulOp_data_0_lpi_1_dfm_mx0_30_0 = cfg_mul_src_1_sva_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10068|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10067" *) chn_mul_op_rsci_d_mxwt[30:0] : cfg_mul_op_1_sva_1[30:0];
  assign FpMul_8U_23U_p_expo_lpi_1_dfm_1_mx0 = FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) FpMul_8U_23U_p_expo_sva_5 : mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  assign FpMul_8U_23U_p_expo_3_lpi_1_dfm_1_mx0 = FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) FpMul_8U_23U_p_expo_3_sva_5 : mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  assign FpMul_8U_23U_p_expo_2_lpi_1_dfm_1_mx0 = FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) FpMul_8U_23U_p_expo_2_sva_5 : mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  assign FpMul_8U_23U_p_expo_1_lpi_1_dfm_1_mx0 = FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10153|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10152" *) FpMul_8U_23U_p_expo_1_sva_5 : mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  assign _00022_ = FpMul_8U_23U_lor_2_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) 23'b11111111111111111111111 : FpMul_8U_23U_nor_6_nl;
  assign _00021_ = _00850_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) mux_240_nl : 23'b11111111111111111111111;
  assign mux_240_nl = or_842_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) mul_mul_4_FpMantRNE_48U_24U_else_acc_nl : { _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22] };
  assign _00019_ = FpMul_8U_23U_lor_11_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) 23'b11111111111111111111111 : FpMul_8U_23U_nor_5_nl;
  assign _00018_ = _00848_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) mux_239_nl : 23'b11111111111111111111111;
  assign mux_239_nl = or_841_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) mul_mul_3_FpMantRNE_48U_24U_else_acc_nl : { _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22] };
  assign _00016_ = FpMul_8U_23U_lor_10_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) 23'b11111111111111111111111 : FpMul_8U_23U_nor_4_nl;
  assign _00015_ = _00846_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) mux_238_nl : 23'b11111111111111111111111;
  assign mux_238_nl = or_840_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) mul_mul_2_FpMantRNE_48U_24U_else_acc_nl : { _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22] };
  assign _00013_ = FpMul_8U_23U_lor_9_lpi_1_dfm ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) 23'b11111111111111111111111 : FpMul_8U_23U_nor_nl;
  assign _00012_ = or_tmp_133 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) mux_237_nl : 23'b11111111111111111111111;
  assign mux_237_nl = or_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10051|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10050" *) mul_mul_1_FpMantRNE_48U_24U_else_acc_nl : { _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22] };
  assign FpMul_8U_23U_p_mant_p1_sva_mx1 = FpMul_8U_23U_p_mant_p1_and_4_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10119|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10118" *) mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp : FpMul_8U_23U_p_mant_p1_sva;
  assign FpMul_8U_23U_p_mant_p1_3_sva_mx1 = FpMul_8U_23U_p_mant_p1_and_5_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10119|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10118" *) mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp : FpMul_8U_23U_p_mant_p1_3_sva;
  assign FpMul_8U_23U_p_mant_p1_2_sva_mx1 = FpMul_8U_23U_p_mant_p1_and_6_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10119|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10118" *) mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp : FpMul_8U_23U_p_mant_p1_2_sva;
  assign FpMul_8U_23U_p_mant_p1_1_sva_mx1 = FpMul_8U_23U_p_mant_p1_and_7_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10119|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10118" *) mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp : FpMul_8U_23U_p_mant_p1_1_sva;
  assign mux_178_nl = and_20_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_496_nl : or_tmp_46;
  assign mux_173_nl = and_20_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_488_nl : or_tmp_29;
  assign mux_168_nl = and_20_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_480_nl : or_tmp_15;
  assign mux_160_nl = and_20_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) or_467_nl : or_tmp_1;
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st : mul_mul_4_FpMantRNE_48U_24U_else_and_tmp;
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st : mul_mul_3_FpMantRNE_48U_24U_else_and_tmp;
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st : mul_mul_2_FpMantRNE_48U_24U_else_and_tmp;
  assign FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st : mul_mul_1_FpMantRNE_48U_24U_else_and_tmp;
  assign mux_33_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_307_nl : nor_308_nl;
  assign mux_31_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_311_nl : nor_312_nl;
  assign mux_29_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_315_nl : nor_316_nl;
  assign mux_27_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) nor_319_nl : nor_320_nl;
  assign mux_26_nl = or_74_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) main_stage_v_2 : main_stage_v_3;
  assign _00277_ = _00608_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9155" *) mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 : mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm;
  assign _00273_ = _00607_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9146" *) mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl[8] : mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  assign _00261_ = _00606_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9136" *) mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 : mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm;
  assign _00257_ = _00605_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9127" *) mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl[8] : mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  assign _00245_ = _00604_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9117" *) mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 : mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm;
  assign _00241_ = _00603_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9108" *) mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl[8] : mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  assign _00229_ = _00602_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9098" *) mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0 : mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm;
  assign _00225_ = _00601_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9089" *) mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl[8] : mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs;
  assign _00172_ = _00600_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9079" *) cfg_mul_src_rsci_d : cfg_mul_src_1_sva_st;
  assign _00143_ = IsNaN_8U_23U_aelse_and_7_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9070" *) IsNaN_8U_23U_land_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_land_lpi_1_dfm_st;
  assign _00164_ = IsNaN_8U_23U_aelse_and_7_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9070" *) IsZero_8U_23U_land_lpi_1_dfm_mx1w0 : IsZero_8U_23U_land_lpi_1_dfm;
  assign _00136_ = IsNaN_8U_23U_aelse_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9060" *) IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_land_3_lpi_1_dfm_st;
  assign _00161_ = IsNaN_8U_23U_aelse_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9060" *) IsZero_8U_23U_land_3_lpi_1_dfm_mx1w0 : IsZero_8U_23U_land_3_lpi_1_dfm;
  assign _00129_ = IsNaN_8U_23U_aelse_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9050" *) IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_land_2_lpi_1_dfm_st;
  assign _00158_ = IsNaN_8U_23U_aelse_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9050" *) IsZero_8U_23U_land_2_lpi_1_dfm_mx1w0 : IsZero_8U_23U_land_2_lpi_1_dfm;
  assign _00122_ = IsNaN_8U_23U_aelse_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9040" *) IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_land_1_lpi_1_dfm_st;
  assign _00155_ = IsNaN_8U_23U_aelse_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9040" *) IsZero_8U_23U_land_1_lpi_1_dfm_mx1w0 : IsZero_8U_23U_land_1_lpi_1_dfm;
  assign _00065_ = _00599_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9031" *) FpMul_8U_23U_lor_1_lpi_1_dfm_mx0w0 : FpMul_8U_23U_lor_1_lpi_1_dfm_st;
  assign _00153_ = _00598_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9023" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp : IsZero_8U_23U_1_land_lpi_1_dfm_5;
  assign _00080_ = _00596_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9015" *) FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0 : FpMul_8U_23U_lor_8_lpi_1_dfm_st;
  assign _00151_ = _00595_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9007" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp : IsZero_8U_23U_1_land_3_lpi_1_dfm_5;
  assign _00075_ = _00593_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8999" *) FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0 : FpMul_8U_23U_lor_7_lpi_1_dfm_st;
  assign _00149_ = _00592_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8991" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp : IsZero_8U_23U_1_land_2_lpi_1_dfm_5;
  assign _00070_ = _00590_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8983" *) FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0 : FpMul_8U_23U_lor_6_lpi_1_dfm_st;
  assign _00147_ = _00589_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8975" *) IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp : IsZero_8U_23U_1_land_1_lpi_1_dfm_5;
  assign _00369_ = and_158_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs : mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign _00274_ = _00587_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8965" *) _00369_ : mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign _00102_ = _00584_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8955" *) mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp : FpMul_8U_23U_p_mant_p1_sva;
  assign _00368_ = and_154_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs : mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign _00258_ = _00582_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8943" *) _00368_ : mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign _00101_ = _00579_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8933" *) mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp : FpMul_8U_23U_p_mant_p1_3_sva;
  assign _00367_ = and_150_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs : mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign _00242_ = _00577_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8922" *) _00367_ : mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign _00100_ = _00574_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8912" *) mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp : FpMul_8U_23U_p_mant_p1_2_sva;
  assign _00175_ = _00572_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8903" *) cfg_truncate_1_sva_1 : cfg_truncate_1_sva_3;
  assign _00366_ = and_146_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs : mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign _00226_ = _00568_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8891" *) _00366_ : mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_2;
  assign _00099_ = _00565_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8881" *) mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp : FpMul_8U_23U_p_mant_p1_1_sva;
  assign _00089_ = _00563_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8869" *) _06024_ : FpMul_8U_23U_mux_49_itm_3;
  assign _00117_ = _00561_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8860" *) IsNaN_8U_23U_1_land_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _00063_ = _00559_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8851" *) _00560_ : FpMul_8U_23U_lor_1_lpi_1_dfm_6;
  assign _00087_ = _00558_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8841" *) _06023_ : FpMul_8U_23U_mux_36_itm_3;
  assign _00115_ = _00556_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8832" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _00078_ = _00554_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8823" *) _00555_ : FpMul_8U_23U_lor_8_lpi_1_dfm_6;
  assign _00085_ = _00553_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8813" *) _06022_ : FpMul_8U_23U_mux_23_itm_3;
  assign _00113_ = _00551_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8804" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _00073_ = _00549_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8795" *) _00550_ : FpMul_8U_23U_lor_7_lpi_1_dfm_6;
  assign _00083_ = _00548_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8785" *) _06021_ : FpMul_8U_23U_mux_10_itm_3;
  assign _00111_ = _00546_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8776" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _00068_ = _00544_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8767" *) _00545_ : FpMul_8U_23U_lor_6_lpi_1_dfm_6;
  assign _00279_ = IntShiftRight_64U_10U_32U_obits_fixed_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8758" *) mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 : mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  assign _00281_ = IntShiftRight_64U_10U_32U_obits_fixed_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8758" *) mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 : mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  assign _00210_ = else_MulOp_data_and_7_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8746" *) else_MulOp_data_3_lpi_1_dfm_2_30_0_1[22:0] : else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm;
  assign _00268_ = else_MulOp_data_and_7_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8746" *) mul_mul_4_FpMantRNE_48U_24U_else_and_tmp : mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st;
  assign _00043_ = else_MulOp_data_and_7_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8746" *) FpMul_8U_23U_FpMul_8U_23U_and_14_itm_mx0w0 : FpMul_8U_23U_FpMul_8U_23U_and_14_itm;
  assign _00037_ = else_MulOp_data_and_7_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8746" *) FpMantRNE_48U_24U_else_carry_sva_mx0w0 : FpMantRNE_48U_24U_else_carry_sva;
  assign _00212_ = _00543_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8735" *) else_MulOp_data_3_lpi_1_dfm_2_30_0_1[30:23] : else_MulOp_data_slc_else_MulOp_data_3_30_23_5_itm;
  assign _00271_ = FpMul_8U_23U_p_expo_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8724" *) mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47] : mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign _00051_ = FpMul_8U_23U_p_expo_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8724" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0 : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm;
  assign _00097_ = FpMul_8U_23U_p_expo_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8724" *) FpMul_8U_23U_p_expo_sva_1_mx0w0 : FpMul_8U_23U_p_expo_sva_1;
  assign _00270_ = _00542_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8713" *) FpMul_8U_23U_p_mant_46_1_lpi_1_dfm_3_mx0[45:23] : mul_mul_4_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  assign _00061_ = _00541_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8703" *) mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] : FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2;
  assign _00263_ = IntShiftRight_64U_10U_32U_obits_fixed_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8693" *) mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 : mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  assign _00265_ = IntShiftRight_64U_10U_32U_obits_fixed_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8693" *) mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 : mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  assign _00207_ = else_MulOp_data_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8681" *) else_MulOp_data_2_lpi_1_dfm_2_30_0_1[22:0] : else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm;
  assign _00252_ = else_MulOp_data_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8681" *) mul_mul_3_FpMantRNE_48U_24U_else_and_tmp : mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st;
  assign _00041_ = else_MulOp_data_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8681" *) FpMul_8U_23U_FpMul_8U_23U_and_13_itm_mx0w0 : FpMul_8U_23U_FpMul_8U_23U_and_13_itm;
  assign _00035_ = else_MulOp_data_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8681" *) FpMantRNE_48U_24U_else_carry_3_sva_mx0w0 : FpMantRNE_48U_24U_else_carry_3_sva;
  assign _00209_ = _00540_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8670" *) else_MulOp_data_2_lpi_1_dfm_2_30_0_1[30:23] : else_MulOp_data_slc_else_MulOp_data_2_30_23_5_itm;
  assign _00255_ = FpMul_8U_23U_p_expo_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8659" *) mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47] : mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign _00049_ = FpMul_8U_23U_p_expo_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8659" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0 : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm;
  assign _00095_ = FpMul_8U_23U_p_expo_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8659" *) FpMul_8U_23U_p_expo_3_sva_1_mx0w0 : FpMul_8U_23U_p_expo_3_sva_1;
  assign _00254_ = _00539_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8648" *) FpMul_8U_23U_p_mant_46_1_3_lpi_1_dfm_3_mx0[45:23] : mul_mul_3_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  assign _00059_ = _00538_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8638" *) mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] : FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2;
  assign _00247_ = IntShiftRight_64U_10U_32U_obits_fixed_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8628" *) mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 : mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  assign _00249_ = IntShiftRight_64U_10U_32U_obits_fixed_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8628" *) mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 : mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  assign _00204_ = else_MulOp_data_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8616" *) else_MulOp_data_1_lpi_1_dfm_2_30_0_1[22:0] : else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm;
  assign _00236_ = else_MulOp_data_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8616" *) mul_mul_2_FpMantRNE_48U_24U_else_and_tmp : mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st;
  assign _00039_ = else_MulOp_data_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8616" *) FpMul_8U_23U_FpMul_8U_23U_and_12_itm_mx0w0 : FpMul_8U_23U_FpMul_8U_23U_and_12_itm;
  assign _00033_ = else_MulOp_data_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8616" *) FpMantRNE_48U_24U_else_carry_2_sva_mx0w0 : FpMantRNE_48U_24U_else_carry_2_sva;
  assign _00206_ = _00537_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8605" *) else_MulOp_data_1_lpi_1_dfm_2_30_0_1[30:23] : else_MulOp_data_slc_else_MulOp_data_1_30_23_5_itm;
  assign _00239_ = FpMul_8U_23U_p_expo_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8594" *) mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47] : mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign _00047_ = FpMul_8U_23U_p_expo_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8594" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0 : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm;
  assign _00093_ = FpMul_8U_23U_p_expo_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8594" *) FpMul_8U_23U_p_expo_2_sva_1_mx0w0 : FpMul_8U_23U_p_expo_2_sva_1;
  assign _00238_ = _00536_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8583" *) FpMul_8U_23U_p_mant_46_1_2_lpi_1_dfm_3_mx0[45:23] : mul_mul_2_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  assign _00057_ = _00535_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8573" *) mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] : FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2;
  assign _00231_ = IntShiftRight_64U_10U_32U_obits_fixed_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8563" *) mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0 : mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm;
  assign _00233_ = IntShiftRight_64U_10U_32U_obits_fixed_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8563" *) mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0 : mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm;
  assign _00201_ = else_MulOp_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8551" *) else_MulOp_data_0_lpi_1_dfm_2_30_0_1[22:0] : else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm;
  assign _00220_ = else_MulOp_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8551" *) mul_mul_1_FpMantRNE_48U_24U_else_and_tmp : mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st;
  assign _00045_ = else_MulOp_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8551" *) FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0 : FpMul_8U_23U_FpMul_8U_23U_and_itm;
  assign _00031_ = else_MulOp_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8551" *) FpMantRNE_48U_24U_else_carry_1_sva_mx0w0 : FpMantRNE_48U_24U_else_carry_1_sva;
  assign _00203_ = _00534_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8540" *) else_MulOp_data_0_lpi_1_dfm_2_30_0_1[30:23] : else_MulOp_data_slc_else_MulOp_data_0_30_23_5_itm;
  assign _00223_ = FpMul_8U_23U_p_expo_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8529" *) mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47] : mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm;
  assign _00053_ = FpMul_8U_23U_p_expo_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8529" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0 : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm;
  assign _00091_ = FpMul_8U_23U_p_expo_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8529" *) FpMul_8U_23U_p_expo_1_sva_1_mx0w0 : FpMul_8U_23U_p_expo_1_sva_1;
  assign _00222_ = _00533_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8518" *) FpMul_8U_23U_p_mant_46_1_1_lpi_1_dfm_3_mx0[45:23] : mul_mul_1_FpMantWidthDec_8U_47U_23U_0U_0U_overflow_slc_FpMantRNE_48U_24U_i_data_46_1_45_23_itm_1;
  assign _00055_ = _00532_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8508" *) mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7] : FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2;
  assign _00365_ = cfg_mul_src_1_sva_st_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) cfg_mul_src_1_sva_st : cfg_mul_src_rsci_d;
  assign _00173_ = _00531_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8498" *) _00365_ : cfg_mul_src_1_sva_st_1;
  assign _00304_ = mul_mul_aelse_and_19_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8486" *) mul_mul_land_lpi_1_dfm_mx1w0 : mul_mul_land_lpi_1_dfm_st_1;
  assign _00298_ = mul_mul_aelse_and_19_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8486" *) mul_mul_land_3_lpi_1_dfm_mx1w0 : mul_mul_land_3_lpi_1_dfm_st_1;
  assign _00292_ = mul_mul_aelse_and_19_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8486" *) mul_mul_land_2_lpi_1_dfm_mx1w0 : mul_mul_land_2_lpi_1_dfm_st_1;
  assign _00286_ = mul_mul_aelse_and_19_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8486" *) mul_mul_land_1_lpi_1_dfm_mx1w0 : mul_mul_land_1_lpi_1_dfm_st_1;
  assign _00364_ = and_dcpl_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsZero_8U_23U_land_lpi_1_dfm : IsZero_8U_23U_land_lpi_1_dfm_mx1w0;
  assign _00363_ = and_dcpl_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsNaN_8U_23U_land_lpi_1_dfm_st : IsNaN_8U_23U_land_lpi_1_dfm_mx0w0;
  assign _00144_ = IsNaN_8U_23U_aelse_and_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8472" *) _00363_ : IsNaN_8U_23U_land_lpi_1_dfm_st_1;
  assign _00165_ = IsNaN_8U_23U_aelse_and_27_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8472" *) _00364_ : IsZero_8U_23U_land_lpi_1_dfm_4;
  assign _00362_ = and_dcpl_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsZero_8U_23U_land_3_lpi_1_dfm : IsZero_8U_23U_land_3_lpi_1_dfm_mx1w0;
  assign _00361_ = and_dcpl_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st : IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0;
  assign _00137_ = IsNaN_8U_23U_aelse_and_26_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8460" *) _00361_ : IsNaN_8U_23U_land_3_lpi_1_dfm_st_1;
  assign _00162_ = IsNaN_8U_23U_aelse_and_26_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8460" *) _00362_ : IsZero_8U_23U_land_3_lpi_1_dfm_4;
  assign _00360_ = and_dcpl_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsZero_8U_23U_land_2_lpi_1_dfm : IsZero_8U_23U_land_2_lpi_1_dfm_mx1w0;
  assign _00359_ = and_dcpl_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st : IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0;
  assign _00130_ = IsNaN_8U_23U_aelse_and_25_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8448" *) _00359_ : IsNaN_8U_23U_land_2_lpi_1_dfm_st_1;
  assign _00159_ = IsNaN_8U_23U_aelse_and_25_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8448" *) _00360_ : IsZero_8U_23U_land_2_lpi_1_dfm_4;
  assign _00171_ = _00529_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8439" *) cfg_mul_src_rsci_d : cfg_mul_src_1_sva_1;
  assign _00170_ = _00528_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8431" *) cfg_mul_op_rsci_d : cfg_mul_op_1_sva_1;
  assign _00358_ = and_dcpl_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsZero_8U_23U_land_1_lpi_1_dfm : IsZero_8U_23U_land_1_lpi_1_dfm_mx1w0;
  assign _00357_ = and_dcpl_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st : IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0;
  assign _00123_ = IsNaN_8U_23U_aelse_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8419" *) _00357_ : IsNaN_8U_23U_land_1_lpi_1_dfm_st_1;
  assign _00156_ = IsNaN_8U_23U_aelse_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8419" *) _00358_ : IsZero_8U_23U_land_1_lpi_1_dfm_4;
  assign _00169_ = MulIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8400" *) chn_mul_in_rsci_d_mxwt : MulIn_data_sva_1;
  assign _00174_ = MulIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8400" *) cfg_truncate_rsci_d : cfg_truncate_1_sva_1;
  assign _00301_ = MulIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8400" *) mul_mul_land_lpi_1_dfm_mx1w0 : mul_mul_land_lpi_1_dfm_2;
  assign _00295_ = MulIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8400" *) mul_mul_land_3_lpi_1_dfm_mx1w0 : mul_mul_land_3_lpi_1_dfm_2;
  assign _00289_ = MulIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8400" *) mul_mul_land_2_lpi_1_dfm_mx1w0 : mul_mul_land_2_lpi_1_dfm_2;
  assign _00283_ = MulIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8400" *) mul_mul_land_1_lpi_1_dfm_mx1w0 : mul_mul_land_1_lpi_1_dfm_2;
  assign _00214_ = MulIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8400" *) cfg_mul_bypass_rsci_d : io_read_cfg_mul_bypass_rsc_svs_st_1;
  assign _00119_ = MulIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8400" *) IsNaN_8U_23U_land_1_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_land_1_lpi_1_dfm_4;
  assign _00126_ = MulIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8400" *) IsNaN_8U_23U_land_2_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_land_2_lpi_1_dfm_4;
  assign _00133_ = MulIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8400" *) IsNaN_8U_23U_land_3_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_land_3_lpi_1_dfm_4;
  assign _00140_ = MulIn_data_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8400" *) IsNaN_8U_23U_land_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_land_lpi_1_dfm_4;
  assign _00216_ = _00527_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8382" *) _00891_ : main_stage_v_1;
  assign _00306_ = mul_mul_aelse_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8371" *) mul_mul_land_lpi_1_dfm_st_4 : mul_mul_land_lpi_1_dfm_st_5;
  assign _00300_ = mul_mul_aelse_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8371" *) mul_mul_land_3_lpi_1_dfm_st_4 : mul_mul_land_3_lpi_1_dfm_st_5;
  assign _00294_ = mul_mul_aelse_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8371" *) mul_mul_land_2_lpi_1_dfm_st_4 : mul_mul_land_2_lpi_1_dfm_st_5;
  assign _00288_ = mul_mul_aelse_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8371" *) mul_mul_land_1_lpi_1_dfm_st_4 : mul_mul_land_1_lpi_1_dfm_st_5;
  assign _00356_ = and_dcpl_52 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm : mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  assign _00355_ = and_dcpl_52 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm : mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  assign _00280_ = IntShiftRight_64U_10U_32U_obits_fixed_and_22_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8357" *) _00355_ : mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign _00282_ = IntShiftRight_64U_10U_32U_obits_fixed_and_22_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8357" *) _00356_ : mul_mul_4_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  assign _00354_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMantRNE_48U_24U_else_carry_sva : FpMantRNE_48U_24U_else_carry_sva_mx0w0;
  assign _00038_ = _00526_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8347" *) _00354_ : FpMantRNE_48U_24U_else_carry_sva_2;
  assign _00269_ = _00525_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8338" *) FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse : mul_mul_4_FpMantRNE_48U_24U_else_and_svs_st_2;
  assign _00064_ = _00524_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8329" *) FpMul_8U_23U_lor_1_lpi_1_dfm_6 : FpMul_8U_23U_lor_1_lpi_1_dfm_7;
  assign _00146_ = IsNaN_8U_23U_aelse_and_23_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8320" *) IsNaN_8U_23U_land_lpi_1_dfm_st_4 : IsNaN_8U_23U_land_lpi_1_dfm_st_5;
  assign _00067_ = IsNaN_8U_23U_aelse_and_23_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8320" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st_3 : FpMul_8U_23U_lor_1_lpi_1_dfm_st_4;
  assign _00211_ = _00523_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8308" *) _06048_ : else_MulOp_data_slc_else_MulOp_data_3_22_0_1_itm_2;
  assign _00353_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_FpMul_8U_23U_and_14_itm : FpMul_8U_23U_FpMul_8U_23U_and_14_itm_mx0w0;
  assign _00044_ = FpMantRNE_48U_24U_else_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8297" *) _00353_ : FpMul_8U_23U_FpMul_8U_23U_and_14_itm_2;
  assign _00267_ = FpMantRNE_48U_24U_else_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8297" *) FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_1_cse : mul_mul_4_FpMantRNE_48U_24U_else_and_svs_2;
  assign _00110_ = IsNaN_8U_23U_1_aelse_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8287" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva[64] : IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_64_1;
  assign _00118_ = IsNaN_8U_23U_1_aelse_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8287" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6 : IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _00276_ = _00522_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8277" *) mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 : mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign _00352_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm : mul_mul_4_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign _00272_ = _00521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8267" *) _00352_ : mul_mul_4_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  assign _00351_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_mx0w0;
  assign _00052_ = _00520_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8257" *) _00351_ : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_3_itm_2;
  assign _00350_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_2 : mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign _00062_ = _00519_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8245" *) _00350_ : FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_sva_st_3;
  assign _00098_ = _00518_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8232" *) _01022_ : FpMul_8U_23U_p_expo_sva_5;
  assign _00349_ = and_dcpl_52 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm : mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  assign _00348_ = and_dcpl_52 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm : mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  assign _00264_ = IntShiftRight_64U_10U_32U_obits_fixed_and_19_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8220" *) _00348_ : mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign _00266_ = IntShiftRight_64U_10U_32U_obits_fixed_and_19_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8220" *) _00349_ : mul_mul_3_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  assign _00347_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMantRNE_48U_24U_else_carry_3_sva : FpMantRNE_48U_24U_else_carry_3_sva_mx0w0;
  assign _00036_ = _00516_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8210" *) _00347_ : FpMantRNE_48U_24U_else_carry_3_sva_2;
  assign _00253_ = _00515_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8201" *) FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse : mul_mul_3_FpMantRNE_48U_24U_else_and_svs_st_2;
  assign _00079_ = _00514_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8192" *) FpMul_8U_23U_lor_8_lpi_1_dfm_6 : FpMul_8U_23U_lor_8_lpi_1_dfm_7;
  assign _00082_ = IsNaN_8U_23U_aelse_and_21_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8183" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st_3 : FpMul_8U_23U_lor_8_lpi_1_dfm_st_4;
  assign _00139_ = IsNaN_8U_23U_aelse_and_21_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8183" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 : IsNaN_8U_23U_land_3_lpi_1_dfm_st_5;
  assign _00208_ = _00513_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8171" *) _06047_ : else_MulOp_data_slc_else_MulOp_data_2_22_0_1_itm_2;
  assign _00346_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_FpMul_8U_23U_and_13_itm : FpMul_8U_23U_FpMul_8U_23U_and_13_itm_mx0w0;
  assign _00042_ = FpMantRNE_48U_24U_else_and_11_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8160" *) _00346_ : FpMul_8U_23U_FpMul_8U_23U_and_13_itm_2;
  assign _00251_ = FpMantRNE_48U_24U_else_and_11_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8160" *) FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_3_cse : mul_mul_3_FpMantRNE_48U_24U_else_and_svs_2;
  assign _00108_ = IsNaN_8U_23U_1_aelse_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8150" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva[64] : IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_64_1;
  assign _00116_ = IsNaN_8U_23U_1_aelse_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8150" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_6 : IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign _00260_ = _00512_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8140" *) mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 : mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign _00345_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm : mul_mul_3_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign _00256_ = _00511_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8130" *) _00345_ : mul_mul_3_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  assign _00344_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_mx0w0;
  assign _00050_ = _00510_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8120" *) _00344_ : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_2_itm_2;
  assign _00343_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_2 : mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign _00060_ = _00509_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8108" *) _00343_ : FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_3_sva_st_3;
  assign _00096_ = _00508_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8095" *) _01021_ : FpMul_8U_23U_p_expo_3_sva_5;
  assign _00342_ = and_dcpl_52 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm : mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  assign _00341_ = and_dcpl_52 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm : mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  assign _00248_ = IntShiftRight_64U_10U_32U_obits_fixed_and_16_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8083" *) _00341_ : mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign _00250_ = IntShiftRight_64U_10U_32U_obits_fixed_and_16_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8083" *) _00342_ : mul_mul_2_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  assign _00340_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMantRNE_48U_24U_else_carry_2_sva : FpMantRNE_48U_24U_else_carry_2_sva_mx0w0;
  assign _00034_ = _00506_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8073" *) _00340_ : FpMantRNE_48U_24U_else_carry_2_sva_2;
  assign _00237_ = _00505_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8064" *) FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse : mul_mul_2_FpMantRNE_48U_24U_else_and_svs_st_2;
  assign _00074_ = _00504_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8055" *) FpMul_8U_23U_lor_7_lpi_1_dfm_6 : FpMul_8U_23U_lor_7_lpi_1_dfm_7;
  assign _00077_ = IsNaN_8U_23U_aelse_and_19_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8046" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st_3 : FpMul_8U_23U_lor_7_lpi_1_dfm_st_4;
  assign _00132_ = IsNaN_8U_23U_aelse_and_19_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8046" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 : IsNaN_8U_23U_land_2_lpi_1_dfm_st_5;
  assign _00205_ = _00503_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8034" *) _06046_ : else_MulOp_data_slc_else_MulOp_data_1_22_0_1_itm_2;
  assign _00339_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_FpMul_8U_23U_and_12_itm : FpMul_8U_23U_FpMul_8U_23U_and_12_itm_mx0w0;
  assign _00040_ = FpMantRNE_48U_24U_else_and_9_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8023" *) _00339_ : FpMul_8U_23U_FpMul_8U_23U_and_12_itm_2;
  assign _00235_ = FpMantRNE_48U_24U_else_and_9_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8023" *) FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_5_cse : mul_mul_2_FpMantRNE_48U_24U_else_and_svs_2;
  assign _00106_ = IsNaN_8U_23U_1_aelse_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8013" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva[64] : IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_64_1;
  assign _00114_ = IsNaN_8U_23U_1_aelse_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8013" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 : IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _00244_ = _00502_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:8003" *) mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 : mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign _00338_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm : mul_mul_2_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign _00240_ = _00501_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7993" *) _00338_ : mul_mul_2_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  assign _00337_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_mx0w0;
  assign _00048_ = _00500_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7983" *) _00337_ : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_1_itm_2;
  assign _00336_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_2 : mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign _00058_ = _00499_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7971" *) _00336_ : FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_2_sva_st_3;
  assign _00094_ = _00498_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7958" *) _01020_ : FpMul_8U_23U_p_expo_2_sva_5;
  assign _00335_ = and_dcpl_52 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm : mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_mx0w0;
  assign _00334_ = and_dcpl_52 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm : mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_mx0w0;
  assign _00232_ = IntShiftRight_64U_10U_32U_obits_fixed_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7946" *) _00334_ : mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nand_itm_2;
  assign _00234_ = IntShiftRight_64U_10U_32U_obits_fixed_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7946" *) _00335_ : mul_mul_1_IntShiftRight_64U_10U_32U_obits_fixed_nor_1_itm_2;
  assign _00333_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMantRNE_48U_24U_else_carry_1_sva : FpMantRNE_48U_24U_else_carry_1_sva_mx0w0;
  assign _00032_ = _00496_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7936" *) _00333_ : FpMantRNE_48U_24U_else_carry_1_sva_2;
  assign _00221_ = _00495_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7927" *) FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse : mul_mul_1_FpMantRNE_48U_24U_else_and_svs_st_2;
  assign _00069_ = _00494_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7918" *) FpMul_8U_23U_lor_6_lpi_1_dfm_6 : FpMul_8U_23U_lor_6_lpi_1_dfm_7;
  assign _00072_ = IsNaN_8U_23U_aelse_and_17_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7909" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st_3 : FpMul_8U_23U_lor_6_lpi_1_dfm_st_4;
  assign _00125_ = IsNaN_8U_23U_aelse_and_17_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7909" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 : IsNaN_8U_23U_land_1_lpi_1_dfm_st_5;
  assign _00202_ = _00493_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7897" *) _06045_ : else_MulOp_data_slc_else_MulOp_data_0_22_0_1_itm_2;
  assign _00332_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_FpMul_8U_23U_and_itm : FpMul_8U_23U_FpMul_8U_23U_and_itm_mx0w0;
  assign _00219_ = FpMantRNE_48U_24U_else_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7886" *) FpMantRNE_48U_24U_else_FpMantRNE_48U_24U_else_mux_7_cse : mul_mul_1_FpMantRNE_48U_24U_else_and_svs_2;
  assign _00046_ = FpMantRNE_48U_24U_else_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7886" *) _00332_ : FpMul_8U_23U_FpMul_8U_23U_and_itm_2;
  assign _00104_ = IsNaN_8U_23U_1_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7876" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva[64] : IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_64_1;
  assign _00112_ = IsNaN_8U_23U_1_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7876" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 : IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign _00228_ = _00492_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7866" *) mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3 : mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_4;
  assign _00331_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm : mul_mul_1_FpMul_8U_23U_p_mant_p1_mul_tmp[47];
  assign _00224_ = _00491_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7856" *) _00331_ : mul_mul_1_FpMul_8U_23U_else_2_else_slc_FpMul_8U_23U_p_mant_p1_47_itm_2;
  assign _00330_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_mx0w0;
  assign _00054_ = _00490_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7846" *) _00330_ : FpMul_8U_23U_else_2_else_FpMul_8U_23U_else_2_else_nand_itm_2;
  assign _00329_ = and_dcpl_47 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_2 : mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign _00056_ = _00489_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7834" *) _00329_ : FpMul_8U_23U_else_2_else_if_if_slc_FpMul_8U_23U_else_2_else_if_if_acc_1_7_mdf_1_sva_st_3;
  assign _00092_ = _00488_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7821" *) _01019_ : FpMul_8U_23U_p_expo_1_sva_5;
  assign _00109_ = IntShiftRight_64U_10U_32U_obits_fixed_and_11_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7811" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva[31:0] : IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva_1_31_0_1;
  assign _00090_ = IntShiftRight_64U_10U_32U_obits_fixed_and_11_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7811" *) FpMul_8U_23U_mux_49_itm_3 : FpMul_8U_23U_mux_49_itm_4;
  assign _00107_ = IntShiftRight_64U_10U_32U_obits_fixed_and_10_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7801" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva[31:0] : IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva_1_31_0_1;
  assign _00088_ = IntShiftRight_64U_10U_32U_obits_fixed_and_10_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7801" *) FpMul_8U_23U_mux_36_itm_3 : FpMul_8U_23U_mux_36_itm_4;
  assign _00105_ = IntShiftRight_64U_10U_32U_obits_fixed_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7791" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva[31:0] : IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva_1_31_0_1;
  assign _00086_ = IntShiftRight_64U_10U_32U_obits_fixed_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7791" *) FpMul_8U_23U_mux_23_itm_3 : FpMul_8U_23U_mux_23_itm_4;
  assign _00103_ = IntShiftRight_64U_10U_32U_obits_fixed_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7781" *) IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva[31:0] : IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva_1_31_0_1;
  assign _00084_ = IntShiftRight_64U_10U_32U_obits_fixed_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7781" *) FpMul_8U_23U_mux_10_itm_3 : FpMul_8U_23U_mux_10_itm_4;
  assign _00168_ = MulIn_data_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7763" *) MulIn_data_sva_132 : MulIn_data_sva_133;
  assign _00303_ = MulIn_data_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7763" *) mul_mul_land_lpi_1_dfm_5 : mul_mul_land_lpi_1_dfm_6;
  assign _00297_ = MulIn_data_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7763" *) mul_mul_land_3_lpi_1_dfm_5 : mul_mul_land_3_lpi_1_dfm_6;
  assign _00291_ = MulIn_data_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7763" *) mul_mul_land_2_lpi_1_dfm_5 : mul_mul_land_2_lpi_1_dfm_6;
  assign _00285_ = MulIn_data_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7763" *) mul_mul_land_1_lpi_1_dfm_5 : mul_mul_land_1_lpi_1_dfm_6;
  assign _00213_ = MulIn_data_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7763" *) io_read_cfg_mul_bypass_rsc_svs_st_4 : io_read_cfg_mul_bypass_rsc_svs_5;
  assign _00121_ = MulIn_data_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7763" *) IsNaN_8U_23U_land_1_lpi_1_dfm_7 : IsNaN_8U_23U_land_1_lpi_1_dfm_8;
  assign _00128_ = MulIn_data_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7763" *) IsNaN_8U_23U_land_2_lpi_1_dfm_7 : IsNaN_8U_23U_land_2_lpi_1_dfm_8;
  assign _00135_ = MulIn_data_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7763" *) IsNaN_8U_23U_land_3_lpi_1_dfm_7 : IsNaN_8U_23U_land_3_lpi_1_dfm_8;
  assign _00142_ = MulIn_data_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7763" *) IsNaN_8U_23U_land_lpi_1_dfm_7 : IsNaN_8U_23U_land_lpi_1_dfm_8;
  assign _00218_ = _00486_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7745" *) _00885_ : main_stage_v_3;
  assign _00305_ = mul_mul_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7734" *) mul_mul_land_lpi_1_dfm_st_1 : mul_mul_land_lpi_1_dfm_st_4;
  assign _00299_ = mul_mul_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7734" *) mul_mul_land_3_lpi_1_dfm_st_1 : mul_mul_land_3_lpi_1_dfm_st_4;
  assign _00293_ = mul_mul_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7734" *) mul_mul_land_2_lpi_1_dfm_st_1 : mul_mul_land_2_lpi_1_dfm_st_4;
  assign _00287_ = mul_mul_aelse_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7734" *) mul_mul_land_1_lpi_1_dfm_st_1 : mul_mul_land_1_lpi_1_dfm_st_4;
  assign _00373_ = and_dcpl_38 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10136|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10135" *) mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm : mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  assign _00328_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_lor_1_lpi_1_dfm_st : FpMul_8U_23U_lor_1_lpi_1_dfm_mx0w0;
  assign _00278_ = FpMul_8U_23U_oelse_1_and_7_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7720" *) _00373_ : mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_2;
  assign _00066_ = FpMul_8U_23U_oelse_1_and_7_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7720" *) _00328_ : FpMul_8U_23U_lor_1_lpi_1_dfm_st_3;
  assign _00327_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs : mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign _00275_ = _00485_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7709" *) _00327_ : mul_mul_4_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign _00200_ = else_MulOp_data_and_11_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7698" *) else_MulOp_data_3_lpi_1_dfm_mx1[30:0] : else_MulOp_data_3_lpi_1_dfm_2_30_0_1;
  assign _00145_ = else_MulOp_data_and_11_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7698" *) IsNaN_8U_23U_land_lpi_1_dfm_st_1 : IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  assign _00326_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsZero_8U_23U_1_land_lpi_1_dfm_5 : IsZero_8U_23U_1_IsZero_8U_23U_1_nor_3_tmp;
  assign _00154_ = _00484_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7688" *) _00326_ : IsZero_8U_23U_1_land_lpi_1_dfm_6;
  assign _00166_ = _00483_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7679" *) IsZero_8U_23U_land_lpi_1_dfm_4 : IsZero_8U_23U_land_lpi_1_dfm_6;
  assign _00372_ = and_dcpl_38 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10136|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10135" *) mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm : mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  assign _00325_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_lor_8_lpi_1_dfm_st : FpMul_8U_23U_lor_8_lpi_1_dfm_mx0w0;
  assign _00081_ = FpMul_8U_23U_oelse_1_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7668" *) _00325_ : FpMul_8U_23U_lor_8_lpi_1_dfm_st_3;
  assign _00262_ = FpMul_8U_23U_oelse_1_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7668" *) _00372_ : mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_2;
  assign _00324_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs : mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign _00259_ = _00482_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7657" *) _00324_ : mul_mul_3_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign _00199_ = else_MulOp_data_and_10_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7646" *) else_MulOp_data_2_lpi_1_dfm_mx1[30:0] : else_MulOp_data_2_lpi_1_dfm_2_30_0_1;
  assign _00138_ = else_MulOp_data_and_10_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7646" *) IsNaN_8U_23U_land_3_lpi_1_dfm_st_1 : IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  assign _00323_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsZero_8U_23U_1_land_3_lpi_1_dfm_5 : IsZero_8U_23U_1_IsZero_8U_23U_1_nor_2_tmp;
  assign _00152_ = _00481_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7636" *) _00323_ : IsZero_8U_23U_1_land_3_lpi_1_dfm_6;
  assign _00163_ = _00480_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7627" *) IsZero_8U_23U_land_3_lpi_1_dfm_4 : IsZero_8U_23U_land_3_lpi_1_dfm_6;
  assign _00371_ = and_dcpl_38 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10136|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10135" *) mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm : mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  assign _00322_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_lor_7_lpi_1_dfm_st : FpMul_8U_23U_lor_7_lpi_1_dfm_mx0w0;
  assign _00076_ = FpMul_8U_23U_oelse_1_and_5_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7616" *) _00322_ : FpMul_8U_23U_lor_7_lpi_1_dfm_st_3;
  assign _00246_ = FpMul_8U_23U_oelse_1_and_5_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7616" *) _00371_ : mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_2;
  assign _00321_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs : mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign _00243_ = _00479_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7605" *) _00321_ : mul_mul_2_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign _00198_ = else_MulOp_data_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7594" *) else_MulOp_data_1_lpi_1_dfm_mx1[30:0] : else_MulOp_data_1_lpi_1_dfm_2_30_0_1;
  assign _00131_ = else_MulOp_data_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7594" *) IsNaN_8U_23U_land_2_lpi_1_dfm_st_1 : IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  assign _00320_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsZero_8U_23U_1_land_2_lpi_1_dfm_5 : IsZero_8U_23U_1_IsZero_8U_23U_1_nor_1_tmp;
  assign _00150_ = _00478_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7584" *) _00320_ : IsZero_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _00160_ = _00477_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7575" *) IsZero_8U_23U_land_2_lpi_1_dfm_4 : IsZero_8U_23U_land_2_lpi_1_dfm_6;
  assign _00370_ = and_dcpl_38 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10136|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10135" *) mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm : mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_mx0w0;
  assign _00319_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) FpMul_8U_23U_lor_6_lpi_1_dfm_st : FpMul_8U_23U_lor_6_lpi_1_dfm_mx0w0;
  assign _00071_ = FpMul_8U_23U_oelse_1_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7564" *) _00319_ : FpMul_8U_23U_lor_6_lpi_1_dfm_st_3;
  assign _00230_ = FpMul_8U_23U_oelse_1_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7564" *) _00370_ : mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_2;
  assign _00318_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs : mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign _00227_ = _00476_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7553" *) _00318_ : mul_mul_1_FpMul_8U_23U_else_2_if_slc_FpMul_8U_23U_else_2_if_acc_8_svs_st_3;
  assign _00197_ = else_MulOp_data_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7542" *) else_MulOp_data_0_lpi_1_dfm_mx1[30:0] : else_MulOp_data_0_lpi_1_dfm_2_30_0_1;
  assign _00124_ = else_MulOp_data_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7542" *) IsNaN_8U_23U_land_1_lpi_1_dfm_st_1 : IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  assign _00317_ = and_dcpl_39 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) IsZero_8U_23U_1_land_1_lpi_1_dfm_5 : IsZero_8U_23U_1_IsZero_8U_23U_1_nor_tmp;
  assign _00148_ = _00475_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7532" *) _00317_ : IsZero_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _00215_ = MulIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7514" *) io_read_cfg_mul_bypass_rsc_svs_st_1 : io_read_cfg_mul_bypass_rsc_svs_st_4;
  assign _00167_ = MulIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7514" *) MulIn_data_sva_1 : MulIn_data_sva_132;
  assign _00120_ = MulIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7514" *) IsNaN_8U_23U_land_1_lpi_1_dfm_4 : IsNaN_8U_23U_land_1_lpi_1_dfm_7;
  assign _00127_ = MulIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7514" *) IsNaN_8U_23U_land_2_lpi_1_dfm_4 : IsNaN_8U_23U_land_2_lpi_1_dfm_7;
  assign _00134_ = MulIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7514" *) IsNaN_8U_23U_land_3_lpi_1_dfm_4 : IsNaN_8U_23U_land_3_lpi_1_dfm_7;
  assign _00141_ = MulIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7514" *) IsNaN_8U_23U_land_lpi_1_dfm_4 : IsNaN_8U_23U_land_lpi_1_dfm_7;
  assign _00302_ = MulIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7514" *) mul_mul_land_lpi_1_dfm_2 : mul_mul_land_lpi_1_dfm_5;
  assign _00296_ = MulIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7514" *) mul_mul_land_3_lpi_1_dfm_2 : mul_mul_land_3_lpi_1_dfm_5;
  assign _00290_ = MulIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7514" *) mul_mul_land_2_lpi_1_dfm_2 : mul_mul_land_2_lpi_1_dfm_5;
  assign _00284_ = MulIn_data_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7514" *) mul_mul_land_1_lpi_1_dfm_2 : mul_mul_land_1_lpi_1_dfm_5;
  assign _00157_ = _00474_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7497" *) IsZero_8U_23U_land_1_lpi_1_dfm_4 : IsZero_8U_23U_land_1_lpi_1_dfm_6;
  assign _00217_ = _00473_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7489" *) _00880_ : main_stage_v_2;
  assign _00179_ = _00472_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7481" *) _00879_ : chn_mul_op_rsci_ld_core_psct;
  assign _00308_ = _00471_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7473" *) _00878_ : reg_chn_mul_out_rsci_ld_core_psct_cse;
  assign _00184_ = chn_mul_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7442" *) _06029_ : chn_mul_out_rsci_d_22_1;
  assign _00185_ = chn_mul_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7442" *) _01015_ : chn_mul_out_rsci_d_30_23;
  assign _00188_ = chn_mul_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7442" *) _06030_ : chn_mul_out_rsci_d_54_33;
  assign _00189_ = chn_mul_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7442" *) _01016_ : chn_mul_out_rsci_d_62_55;
  assign _00192_ = chn_mul_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7442" *) _06031_ : chn_mul_out_rsci_d_86_65;
  assign _00193_ = chn_mul_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7442" *) _01017_ : chn_mul_out_rsci_d_94_87;
  assign _00181_ = chn_mul_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7442" *) _06032_ : chn_mul_out_rsci_d_118_97;
  assign _00182_ = chn_mul_out_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7442" *) _01018_ : chn_mul_out_rsci_d_126_119;
  assign _00316_ = and_dcpl_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_mux_115_nl : MulIn_data_sva_133[127];
  assign _00315_ = and_dcpl_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_mux_114_nl : MulIn_data_sva_133[96];
  assign _00314_ = and_dcpl_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_mux_113_nl : MulIn_data_sva_133[95];
  assign _00313_ = and_dcpl_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_mux_112_nl : MulIn_data_sva_133[64];
  assign _00312_ = and_dcpl_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_mux_111_nl : MulIn_data_sva_133[63];
  assign _00311_ = and_dcpl_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_mux_110_nl : MulIn_data_sva_133[32];
  assign _00310_ = and_dcpl_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_mux_109_nl : MulIn_data_sva_133[31];
  assign _00309_ = and_dcpl_22 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10017|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:10016" *) mul_mul_mux_108_nl : MulIn_data_sva_133[0];
  assign _00180_ = chn_mul_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7412" *) _00309_ : chn_mul_out_rsci_d_0;
  assign _00186_ = chn_mul_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7412" *) _00310_ : chn_mul_out_rsci_d_31;
  assign _00187_ = chn_mul_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7412" *) _00311_ : chn_mul_out_rsci_d_32;
  assign _00190_ = chn_mul_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7412" *) _00312_ : chn_mul_out_rsci_d_63;
  assign _00191_ = chn_mul_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7412" *) _00313_ : chn_mul_out_rsci_d_64;
  assign _00194_ = chn_mul_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7412" *) _00314_ : chn_mul_out_rsci_d_95;
  assign _00195_ = chn_mul_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7412" *) _00315_ : chn_mul_out_rsci_d_96;
  assign _00183_ = chn_mul_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7412" *) _00316_ : chn_mul_out_rsci_d_127;
  assign _00177_ = _00470_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7397" *) chn_mul_in_rsci_ld_core_psct_mx0c0 : chn_mul_in_rsci_ld_core_psct;
  assign _00307_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7386" *) or_tmp_587 : reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse;
  assign _00176_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7386" *) _00877_ : chn_mul_in_rsci_iswt0;
  assign _00178_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7386" *) or_tmp_588 : chn_mul_op_rsci_iswt0;
  assign _00196_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:7386" *) and_dcpl_24 : chn_mul_out_rsci_iswt0;
  assign mul_mul_1_FpMul_8U_23U_xor_nl = MulIn_data_sva_1[31] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9822" *) else_MulOp_data_0_lpi_1_dfm_mx1[31];
  assign mul_mul_2_FpMul_8U_23U_xor_nl = MulIn_data_sva_1[63] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9840" *) else_MulOp_data_1_lpi_1_dfm_mx1[31];
  assign mul_mul_3_FpMul_8U_23U_xor_nl = MulIn_data_sva_1[95] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9858" *) else_MulOp_data_2_lpi_1_dfm_mx1[31];
  assign mul_mul_4_FpMul_8U_23U_xor_nl = MulIn_data_sva_1[127] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:9876" *) else_MulOp_data_3_lpi_1_dfm_mx1[31];
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4241" *)
  SDP_Y_CORE_Y_mul_core_cfg_mul_bypass_rsc_triosy_obj Y_mul_core_cfg_mul_bypass_rsc_triosy_obj_inst (
    .cfg_mul_bypass_rsc_triosy_lz(cfg_mul_bypass_rsc_triosy_lz),
    .cfg_mul_bypass_rsc_triosy_obj_bawt(cfg_mul_bypass_rsc_triosy_obj_bawt),
    .cfg_mul_bypass_rsc_triosy_obj_iswt0(reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse),
    .cfg_mul_bypass_rsc_triosy_obj_oswt(cfg_mul_bypass_rsc_triosy_obj_oswt),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4274" *)
  SDP_Y_CORE_Y_mul_core_cfg_mul_op_rsc_triosy_obj Y_mul_core_cfg_mul_op_rsc_triosy_obj_inst (
    .cfg_mul_op_rsc_triosy_lz(cfg_mul_op_rsc_triosy_lz),
    .cfg_mul_op_rsc_triosy_obj_bawt(cfg_mul_op_rsc_triosy_obj_bawt),
    .cfg_mul_op_rsc_triosy_obj_iswt0(reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse),
    .cfg_mul_op_rsc_triosy_obj_oswt(cfg_mul_op_rsc_triosy_obj_oswt),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4252" *)
  SDP_Y_CORE_Y_mul_core_cfg_mul_prelu_rsc_triosy_obj Y_mul_core_cfg_mul_prelu_rsc_triosy_obj_inst (
    .cfg_mul_prelu_rsc_triosy_lz(cfg_mul_prelu_rsc_triosy_lz),
    .cfg_mul_prelu_rsc_triosy_obj_bawt(cfg_mul_prelu_rsc_triosy_obj_bawt),
    .cfg_mul_prelu_rsc_triosy_obj_iswt0(reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse),
    .cfg_mul_prelu_rsc_triosy_obj_oswt(cfg_mul_prelu_rsc_triosy_obj_oswt),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4263" *)
  SDP_Y_CORE_Y_mul_core_cfg_mul_src_rsc_triosy_obj Y_mul_core_cfg_mul_src_rsc_triosy_obj_inst (
    .cfg_mul_src_rsc_triosy_lz(cfg_mul_src_rsc_triosy_lz),
    .cfg_mul_src_rsc_triosy_obj_bawt(cfg_mul_src_rsc_triosy_obj_bawt),
    .cfg_mul_src_rsc_triosy_obj_iswt0(reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse),
    .cfg_mul_src_rsc_triosy_obj_oswt(cfg_mul_src_rsc_triosy_obj_oswt),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4285" *)
  SDP_Y_CORE_Y_mul_core_cfg_truncate_rsc_triosy_obj Y_mul_core_cfg_truncate_rsc_triosy_obj_inst (
    .cfg_truncate_rsc_triosy_lz(cfg_truncate_rsc_triosy_lz),
    .cfg_truncate_rsc_triosy_obj_bawt(cfg_truncate_rsc_triosy_obj_bawt),
    .cfg_truncate_rsc_triosy_obj_iswt0(reg_cfg_truncate_rsc_triosy_obj_ld_core_psct_cse),
    .cfg_truncate_rsc_triosy_obj_oswt(cfg_truncate_rsc_triosy_obj_oswt),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4196" *)
  SDP_Y_CORE_Y_mul_core_chn_mul_in_rsci Y_mul_core_chn_mul_in_rsci_inst (
    .chn_mul_in_rsc_lz(chn_mul_in_rsc_lz),
    .chn_mul_in_rsc_vz(chn_mul_in_rsc_vz),
    .chn_mul_in_rsc_z(chn_mul_in_rsc_z),
    .chn_mul_in_rsci_bawt(chn_mul_in_rsci_bawt),
    .chn_mul_in_rsci_d_mxwt(chn_mul_in_rsci_d_mxwt),
    .chn_mul_in_rsci_iswt0(chn_mul_in_rsci_iswt0),
    .chn_mul_in_rsci_ld_core_psct(chn_mul_in_rsci_ld_core_psct),
    .chn_mul_in_rsci_oswt(chn_mul_in_rsci_oswt),
    .chn_mul_in_rsci_wen_comp(chn_mul_in_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4211" *)
  SDP_Y_CORE_Y_mul_core_chn_mul_op_rsci Y_mul_core_chn_mul_op_rsci_inst (
    .chn_mul_op_rsc_lz(chn_mul_op_rsc_lz),
    .chn_mul_op_rsc_vz(chn_mul_op_rsc_vz),
    .chn_mul_op_rsc_z(chn_mul_op_rsc_z),
    .chn_mul_op_rsci_bawt(chn_mul_op_rsci_bawt),
    .chn_mul_op_rsci_d_mxwt(chn_mul_op_rsci_d_mxwt),
    .chn_mul_op_rsci_iswt0(chn_mul_op_rsci_iswt0),
    .chn_mul_op_rsci_ld_core_psct(chn_mul_op_rsci_ld_core_psct),
    .chn_mul_op_rsci_oswt(chn_mul_op_rsci_oswt),
    .chn_mul_op_rsci_wen_comp(chn_mul_op_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4226" *)
  SDP_Y_CORE_Y_mul_core_chn_mul_out_rsci Y_mul_core_chn_mul_out_rsci_inst (
    .chn_mul_out_rsc_lz(chn_mul_out_rsc_lz),
    .chn_mul_out_rsc_vz(chn_mul_out_rsc_vz),
    .chn_mul_out_rsc_z(chn_mul_out_rsc_z),
    .chn_mul_out_rsci_bawt(chn_mul_out_rsci_bawt),
    .chn_mul_out_rsci_d({ chn_mul_out_rsci_d_127, chn_mul_out_rsci_d_126_119, chn_mul_out_rsci_d_118_97, chn_mul_out_rsci_d_96, chn_mul_out_rsci_d_95, chn_mul_out_rsci_d_94_87, chn_mul_out_rsci_d_86_65, chn_mul_out_rsci_d_64, chn_mul_out_rsci_d_63, chn_mul_out_rsci_d_62_55, chn_mul_out_rsci_d_54_33, chn_mul_out_rsci_d_32, chn_mul_out_rsci_d_31, chn_mul_out_rsci_d_30_23, chn_mul_out_rsci_d_22_1, chn_mul_out_rsci_d_0 }),
    .chn_mul_out_rsci_iswt0(chn_mul_out_rsci_iswt0),
    .chn_mul_out_rsci_ld_core_psct(reg_chn_mul_out_rsci_ld_core_psct_cse),
    .chn_mul_out_rsci_oswt(chn_mul_out_rsci_oswt),
    .chn_mul_out_rsci_wen_comp(chn_mul_out_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4305" *)
  SDP_Y_CORE_Y_mul_core_core_fsm Y_mul_core_core_fsm_inst (
    .core_wen(core_wen),
    .fsm_output(fsm_output),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4296" *)
  SDP_Y_CORE_Y_mul_core_staller Y_mul_core_staller_inst (
    .chn_mul_in_rsci_wen_comp(chn_mul_in_rsci_wen_comp),
    .chn_mul_op_rsci_wen_comp(chn_mul_op_rsci_wen_comp),
    .chn_mul_out_rsci_wen_comp(chn_mul_out_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4160" *)
  \$paramod\SDP_Y_CORE_mgc_shift_r_v4\width_a=1087\signd_a=1\width_s=10\width_z=1087  mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg (
    .a({ mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_2, 1023'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_3),
    .z(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4169" *)
  \$paramod\SDP_Y_CORE_mgc_shift_r_v4\width_a=1087\signd_a=1\width_s=10\width_z=1087  mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg (
    .a({ mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_2, 1023'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_3),
    .z(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_2_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4178" *)
  \$paramod\SDP_Y_CORE_mgc_shift_r_v4\width_a=1087\signd_a=1\width_s=10\width_z=1087  mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg (
    .a({ mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_2, 1023'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_3),
    .z(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_3_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:4187" *)
  \$paramod\SDP_Y_CORE_mgc_shift_r_v4\width_a=1087\signd_a=1\width_s=10\width_z=1087  mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg (
    .a({ mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_2, 1023'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_truncate_1_sva_3),
    .z(IntShiftRight_64U_10U_32U_obits_fixed_asn_rndi_sva)
  );
  assign _00011_[21:0] = { _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22], _00011_[22] };
  assign _00014_[21:0] = { _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22], _00014_[22] };
  assign _00017_[21:0] = { _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22], _00017_[22] };
  assign _00020_[21:0] = { _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22], _00020_[22] };
  assign cfg_mul_bypass_rsc_triosy_obj_oswt_unreg_pff = or_tmp_591;
  assign chn_mul_in_rsci_oswt_unreg = or_tmp_587;
  assign chn_mul_op_rsci_oswt_unreg = and_dcpl_30;
  assign mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1 = mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign mul_mul_1_FpMul_8U_23U_else_2_if_acc_itm_8_1 = mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign mul_mul_1_FpMul_8U_23U_oelse_1_acc_itm_9_1 = mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1 = mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign mul_mul_2_FpMul_8U_23U_else_2_if_acc_itm_8_1 = mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign mul_mul_2_FpMul_8U_23U_oelse_1_acc_itm_9_1 = mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1 = mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign mul_mul_3_FpMul_8U_23U_else_2_if_acc_itm_8_1 = mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign mul_mul_3_FpMul_8U_23U_oelse_1_acc_itm_9_1 = mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_itm_7_1 = mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7];
  assign mul_mul_4_FpMul_8U_23U_else_2_if_acc_itm_8_1 = mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl[8];
  assign mul_mul_4_FpMul_8U_23U_oelse_1_acc_itm_9_1 = mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl[9];
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1[7:0] = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_1_sva_1;
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1[7:0] = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_2_sva_1;
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1[7:0] = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_3_sva_1;
  assign nl_FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1[7:0] = FpMantWidthDec_8U_47U_23U_0U_0U_o_expo_sva_1;
  assign nl_FpMul_8U_23U_else_2_else_acc_2_nl[7:0] = FpMul_8U_23U_else_2_else_acc_2_nl;
  assign nl_FpMul_8U_23U_else_2_else_acc_3_nl[7:0] = FpMul_8U_23U_else_2_else_acc_3_nl;
  assign nl_FpMul_8U_23U_else_2_else_acc_4_nl[7:0] = FpMul_8U_23U_else_2_else_acc_4_nl;
  assign nl_FpMul_8U_23U_else_2_else_acc_nl[7:0] = FpMul_8U_23U_else_2_else_acc_nl;
  assign nl_FpMul_8U_23U_oelse_1_acc_1_nl[8:0] = FpMul_8U_23U_oelse_1_acc_1_nl;
  assign nl_FpMul_8U_23U_oelse_1_acc_2_nl[8:0] = FpMul_8U_23U_oelse_1_acc_2_nl;
  assign nl_FpMul_8U_23U_oelse_1_acc_3_nl[8:0] = FpMul_8U_23U_oelse_1_acc_3_nl;
  assign nl_FpMul_8U_23U_oelse_1_acc_nl[8:0] = FpMul_8U_23U_oelse_1_acc_nl;
  assign nl_FpMul_8U_23U_p_expo_1_sva_1_mx0w0[7:0] = FpMul_8U_23U_p_expo_1_sva_1_mx0w0;
  assign nl_FpMul_8U_23U_p_expo_2_sva_1_mx0w0[7:0] = FpMul_8U_23U_p_expo_2_sva_1_mx0w0;
  assign nl_FpMul_8U_23U_p_expo_3_sva_1_mx0w0[7:0] = FpMul_8U_23U_p_expo_3_sva_1_mx0w0;
  assign nl_FpMul_8U_23U_p_expo_sva_1_mx0w0[7:0] = FpMul_8U_23U_p_expo_sva_1_mx0w0;
  assign nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva[64:0] = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_1_sva;
  assign nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva[64:0] = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_2_sva;
  assign nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva[64:0] = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_3_sva;
  assign nl_IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva[64:0] = IntShiftRight_64U_10U_32U_obits_fixed_acc_sat_sva;
  assign nl_Y_mul_core_chn_mul_out_rsci_inst_chn_mul_out_rsci_d = { chn_mul_out_rsci_d_127, chn_mul_out_rsci_d_126_119, chn_mul_out_rsci_d_118_97, chn_mul_out_rsci_d_96, chn_mul_out_rsci_d_95, chn_mul_out_rsci_d_94_87, chn_mul_out_rsci_d_86_65, chn_mul_out_rsci_d_64, chn_mul_out_rsci_d_63, chn_mul_out_rsci_d_62_55, chn_mul_out_rsci_d_54_33, chn_mul_out_rsci_d_32, chn_mul_out_rsci_d_31, chn_mul_out_rsci_d_30_23, chn_mul_out_rsci_d_22_1, chn_mul_out_rsci_d_0 };
  assign nl_mul_mul_1_FpMantRNE_48U_24U_else_acc_nl[22:0] = mul_mul_1_FpMantRNE_48U_24U_else_acc_nl;
  assign nl_mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl[8:0] = mul_mul_1_FpMul_8U_23U_else_2_acc_1_nl;
  assign nl_mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0] = mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  assign nl_mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0] = mul_mul_1_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  assign nl_mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl[8:0] = mul_mul_1_FpMul_8U_23U_else_2_if_acc_nl;
  assign nl_mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl[9:0] = mul_mul_1_FpMul_8U_23U_oelse_1_acc_nl;
  assign nl_mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a = { mul_mul_1_IntMulExt_32U_32U_64U_o_mul_itm_2, 1023'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_mul_mul_1_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s = cfg_truncate_1_sva_3;
  assign nl_mul_mul_2_FpMantRNE_48U_24U_else_acc_nl[22:0] = mul_mul_2_FpMantRNE_48U_24U_else_acc_nl;
  assign nl_mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl[8:0] = mul_mul_2_FpMul_8U_23U_else_2_acc_1_nl;
  assign nl_mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0] = mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  assign nl_mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0] = mul_mul_2_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  assign nl_mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl[8:0] = mul_mul_2_FpMul_8U_23U_else_2_if_acc_nl;
  assign nl_mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl[9:0] = mul_mul_2_FpMul_8U_23U_oelse_1_acc_nl;
  assign nl_mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a = { mul_mul_2_IntMulExt_32U_32U_64U_o_mul_itm_2, 1023'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_mul_mul_2_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s = cfg_truncate_1_sva_3;
  assign nl_mul_mul_3_FpMantRNE_48U_24U_else_acc_nl[22:0] = mul_mul_3_FpMantRNE_48U_24U_else_acc_nl;
  assign nl_mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl[8:0] = mul_mul_3_FpMul_8U_23U_else_2_acc_1_nl;
  assign nl_mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0] = mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  assign nl_mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0] = mul_mul_3_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  assign nl_mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl[8:0] = mul_mul_3_FpMul_8U_23U_else_2_if_acc_nl;
  assign nl_mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl[9:0] = mul_mul_3_FpMul_8U_23U_oelse_1_acc_nl;
  assign nl_mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a = { mul_mul_3_IntMulExt_32U_32U_64U_o_mul_itm_2, 1023'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_mul_mul_3_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s = cfg_truncate_1_sva_3;
  assign nl_mul_mul_4_FpMantRNE_48U_24U_else_acc_nl[22:0] = mul_mul_4_FpMantRNE_48U_24U_else_acc_nl;
  assign nl_mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl[8:0] = mul_mul_4_FpMul_8U_23U_else_2_acc_1_nl;
  assign nl_mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl[7:0] = mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_1_nl;
  assign nl_mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl[7:0] = mul_mul_4_FpMul_8U_23U_else_2_else_if_if_acc_nl;
  assign nl_mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl[8:0] = mul_mul_4_FpMul_8U_23U_else_2_if_acc_nl;
  assign nl_mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl[9:0] = mul_mul_4_FpMul_8U_23U_oelse_1_acc_nl;
  assign nl_mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_a = { mul_mul_4_IntMulExt_32U_32U_64U_o_mul_itm_2, 1023'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_mul_mul_4_IntShiftRight_64U_10U_32U_mbits_fixed_rshift_rg_s = cfg_truncate_1_sva_3;
endmodule
