module FP17_ADD_chn_b_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp17_add.v:288" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:289" *)
  output outsig;
  assign outsig = in_0;
endmodule
