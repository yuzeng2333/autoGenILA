module \$paramod\FP17_TO_FP16_mgc_out_stdreg_wait_v1\rscid=2\width=16 (ld, vd, d, lz, vz, z);
  (* src = "./vmod/vlibs/HLS_fp17_to_fp16.v:47" *)
  input [15:0] d;
  (* src = "./vmod/vlibs/HLS_fp17_to_fp16.v:45" *)
  input ld;
  (* src = "./vmod/vlibs/HLS_fp17_to_fp16.v:48" *)
  output lz;
  (* src = "./vmod/vlibs/HLS_fp17_to_fp16.v:46" *)
  output vd;
  (* src = "./vmod/vlibs/HLS_fp17_to_fp16.v:49" *)
  input vz;
  (* src = "./vmod/vlibs/HLS_fp17_to_fp16.v:50" *)
  output [15:0] z;
  assign lz = ld;
  assign vd = vz;
  assign z = d;
endmodule
