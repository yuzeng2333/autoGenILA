module \$paramod\SDP_C_mgc_in_wire_v1\rscid=3\width=16 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:78" *)
  output [15:0] d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:79" *)
  input [15:0] z;
  assign d = z;
endmodule
