module \$paramod\CDP_ICVT_mgc_in_wire_v1\rscid=3\width=16 (d, z);
  (* src = "./vmod/vlibs/HLS_cdp_icvt.v:78" *)
  output [15:0] d;
  (* src = "./vmod/vlibs/HLS_cdp_icvt.v:79" *)
  input [15:0] z;
  assign d = z;
endmodule
