module \$paramod\CDP_OCVT_mgc_in_wire_v1\rscid=2\width=32 (d, z);
  (* src = "./vmod/vlibs/HLS_cdp_ocvt.v:78" *)
  output [31:0] d;
  (* src = "./vmod/vlibs/HLS_cdp_ocvt.v:79" *)
  input [31:0] z;
  assign d = z;
endmodule
