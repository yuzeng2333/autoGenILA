module FP32_TO_FP17_chn_a_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp32_to_fp17.v:166" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp32_to_fp17.v:167" *)
  output outsig;
  assign outsig = in_0;
endmodule
