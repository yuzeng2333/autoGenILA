module ShiftRegister(clock, io_input, io_enable, io_rev, io_cyc, io_tap, io_output_0, io_output_1, io_output_2, io_output_3, io_output_4, io_output_5, io_output_6, io_output_7, io_output_8, io_output_9, io_output_10, io_output_11, io_output_12, io_output_13, io_output_14);
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _000_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _001_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _002_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _003_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _004_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _005_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _006_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _007_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _008_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _009_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _010_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _011_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _012_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _013_;
  (* src = "crypto_accelerator.v:160" *)
  wire [127:0] _014_;
  (* src = "crypto_accelerator.v:165" *)
  wire _015_;
  (* src = "crypto_accelerator.v:176" *)
  wire _016_;
  (* src = "crypto_accelerator.v:189" *)
  wire _017_;
  (* src = "crypto_accelerator.v:202" *)
  wire _018_;
  (* src = "crypto_accelerator.v:215" *)
  wire _019_;
  (* src = "crypto_accelerator.v:228" *)
  wire _020_;
  (* src = "crypto_accelerator.v:241" *)
  wire _021_;
  (* src = "crypto_accelerator.v:254" *)
  wire _022_;
  wire [127:0] _023_;
  wire [127:0] _024_;
  wire [127:0] _025_;
  wire [127:0] _026_;
  wire [127:0] _027_;
  wire [127:0] _028_;
  wire [127:0] _029_;
  wire [127:0] _030_;
  wire [127:0] _031_;
  wire [127:0] _032_;
  wire [127:0] _033_;
  wire [127:0] _034_;
  wire [127:0] _035_;
  wire [127:0] _036_;
  wire [127:0] _037_;
  wire [127:0] _038_;
  wire [127:0] _039_;
  wire [127:0] _040_;
  wire [127:0] _041_;
  wire [127:0] _042_;
  wire [127:0] _043_;
  wire [127:0] _044_;
  wire [127:0] _045_;
  wire [127:0] _046_;
  wire [127:0] _047_;
  wire [127:0] _048_;
  wire [127:0] _049_;
  wire [127:0] _050_;
  wire [127:0] _051_;
  wire [127:0] _052_;
  wire [127:0] _053_;
  wire [127:0] _054_;
  wire [127:0] _055_;
  wire [127:0] _056_;
  wire [127:0] _057_;
  wire [127:0] _058_;
  wire [127:0] _059_;
  wire [127:0] _060_;
  (* src = "crypto_accelerator.v:72" *)
  wire [3:0] _GEN_75;
  (* src = "crypto_accelerator.v:71" *)
  wire [2:0] _T;
  (* src = "crypto_accelerator.v:17" *)
  input clock;
  (* src = "crypto_accelerator.v:21" *)
  input io_cyc;
  (* src = "crypto_accelerator.v:19" *)
  input io_enable;
  (* src = "crypto_accelerator.v:18" *)
  input [127:0] io_input;
  (* src = "crypto_accelerator.v:23" *)
  output [127:0] io_output_0;
  (* src = "crypto_accelerator.v:24" *)
  output [127:0] io_output_1;
  (* src = "crypto_accelerator.v:33" *)
  output [127:0] io_output_10;
  (* src = "crypto_accelerator.v:34" *)
  output [127:0] io_output_11;
  (* src = "crypto_accelerator.v:35" *)
  output [127:0] io_output_12;
  (* src = "crypto_accelerator.v:36" *)
  output [127:0] io_output_13;
  (* src = "crypto_accelerator.v:37" *)
  output [127:0] io_output_14;
  (* src = "crypto_accelerator.v:25" *)
  output [127:0] io_output_2;
  (* src = "crypto_accelerator.v:26" *)
  output [127:0] io_output_3;
  (* src = "crypto_accelerator.v:27" *)
  output [127:0] io_output_4;
  (* src = "crypto_accelerator.v:28" *)
  output [127:0] io_output_5;
  (* src = "crypto_accelerator.v:29" *)
  output [127:0] io_output_6;
  (* src = "crypto_accelerator.v:30" *)
  output [127:0] io_output_7;
  (* src = "crypto_accelerator.v:31" *)
  output [127:0] io_output_8;
  (* src = "crypto_accelerator.v:32" *)
  output [127:0] io_output_9;
  (* src = "crypto_accelerator.v:20" *)
  input io_rev;
  (* src = "crypto_accelerator.v:22" *)
  input io_tap;
  (* src = "crypto_accelerator.v:56" *)
  reg [127:0] reg_0;
  (* src = "crypto_accelerator.v:57" *)
  reg [127:0] reg_1;
  (* src = "crypto_accelerator.v:66" *)
  reg [127:0] reg_10;
  (* src = "crypto_accelerator.v:67" *)
  reg [127:0] reg_11;
  (* src = "crypto_accelerator.v:68" *)
  reg [127:0] reg_12;
  (* src = "crypto_accelerator.v:69" *)
  reg [127:0] reg_13;
  (* src = "crypto_accelerator.v:70" *)
  reg [127:0] reg_14;
  (* src = "crypto_accelerator.v:58" *)
  reg [127:0] reg_2;
  (* src = "crypto_accelerator.v:59" *)
  reg [127:0] reg_3;
  (* src = "crypto_accelerator.v:60" *)
  reg [127:0] reg_4;
  (* src = "crypto_accelerator.v:61" *)
  reg [127:0] reg_5;
  (* src = "crypto_accelerator.v:62" *)
  reg [127:0] reg_6;
  (* src = "crypto_accelerator.v:63" *)
  reg [127:0] reg_7;
  (* src = "crypto_accelerator.v:64" *)
  reg [127:0] reg_8;
  (* src = "crypto_accelerator.v:65" *)
  reg [127:0] reg_9;
  assign _015_ = ! (* src = "crypto_accelerator.v:165" *) _T;
  assign _016_ = 1'b1 == (* src = "crypto_accelerator.v:176" *) _T;
  assign _017_ = 2'b10 == (* src = "crypto_accelerator.v:189" *) _T;
  assign _018_ = 2'b11 == (* src = "crypto_accelerator.v:202" *) _T;
  assign _019_ = 3'b100 == (* src = "crypto_accelerator.v:215" *) _T;
  assign _021_ = 3'b110 == (* src = "crypto_accelerator.v:241" *) _T;
  assign _022_ = 3'b111 == (* src = "crypto_accelerator.v:254" *) _T;
  assign _020_ = 3'b101 == (* src = "crypto_accelerator.v:360" *) _T;
  always @(posedge clock)
      reg_0 <= _000_;
  always @(posedge clock)
      reg_1 <= _006_;
  always @(posedge clock)
      reg_2 <= _007_;
  always @(posedge clock)
      reg_3 <= _008_;
  always @(posedge clock)
      reg_4 <= _009_;
  always @(posedge clock)
      reg_5 <= _010_;
  always @(posedge clock)
      reg_6 <= _011_;
  always @(posedge clock)
      reg_7 <= _012_;
  always @(posedge clock)
      reg_8 <= _013_;
  always @(posedge clock)
      reg_9 <= _014_;
  always @(posedge clock)
      reg_10 <= _001_;
  always @(posedge clock)
      reg_11 <= _002_;
  always @(posedge clock)
      reg_12 <= _003_;
  always @(posedge clock)
      reg_13 <= _004_;
  always @(posedge clock)
      reg_14 <= _005_;
  assign _023_ = _016_ ? (* src = "crypto_accelerator.v:368" *) reg_1 : reg_0;
  assign _024_ = _017_ ? (* src = "crypto_accelerator.v:366" *) reg_2 : _023_;
  assign _025_ = _018_ ? (* src = "crypto_accelerator.v:364" *) reg_3 : _024_;
  assign _026_ = _019_ ? (* src = "crypto_accelerator.v:362" *) reg_4 : _025_;
  assign _027_ = _020_ ? (* src = "crypto_accelerator.v:360" *) reg_5 : _026_;
  assign _028_ = _021_ ? (* src = "crypto_accelerator.v:358" *) reg_6 : _027_;
  assign _029_ = _022_ ? (* src = "crypto_accelerator.v:356" *) reg_7 : _028_;
  assign _030_ = io_rev ? (* src = "crypto_accelerator.v:342" *) _029_ : reg_13;
  assign _005_ = io_enable ? (* src = "crypto_accelerator.v:341" *) _030_ : reg_14;
  assign _031_ = io_rev ? (* src = "crypto_accelerator.v:329" *) reg_14 : reg_12;
  assign _004_ = io_enable ? (* src = "crypto_accelerator.v:328" *) _031_ : reg_13;
  assign _032_ = io_rev ? (* src = "crypto_accelerator.v:316" *) reg_13 : reg_11;
  assign _003_ = io_enable ? (* src = "crypto_accelerator.v:315" *) _032_ : reg_12;
  assign _033_ = io_rev ? (* src = "crypto_accelerator.v:303" *) reg_12 : reg_10;
  assign _002_ = io_enable ? (* src = "crypto_accelerator.v:302" *) _033_ : reg_11;
  assign _034_ = io_rev ? (* src = "crypto_accelerator.v:290" *) reg_11 : reg_9;
  assign _001_ = io_enable ? (* src = "crypto_accelerator.v:289" *) _034_ : reg_10;
  assign _035_ = io_rev ? (* src = "crypto_accelerator.v:277" *) reg_10 : reg_8;
  assign _014_ = io_enable ? (* src = "crypto_accelerator.v:276" *) _035_ : reg_9;
  assign _036_ = io_rev ? (* src = "crypto_accelerator.v:264" *) reg_9 : reg_7;
  assign _013_ = io_enable ? (* src = "crypto_accelerator.v:263" *) _036_ : reg_8;
  assign _037_ = _022_ ? (* src = "crypto_accelerator.v:254" *) reg_14 : reg_6;
  assign _038_ = io_cyc ? (* src = "crypto_accelerator.v:253" *) _037_ : reg_6;
  assign _039_ = io_rev ? (* src = "crypto_accelerator.v:251" *) reg_8 : _038_;
  assign _012_ = io_enable ? (* src = "crypto_accelerator.v:250" *) _039_ : reg_7;
  assign _040_ = _021_ ? (* src = "crypto_accelerator.v:241" *) reg_14 : reg_5;
  assign _041_ = io_cyc ? (* src = "crypto_accelerator.v:240" *) _040_ : reg_5;
  assign _042_ = io_rev ? (* src = "crypto_accelerator.v:238" *) reg_7 : _041_;
  assign _011_ = io_enable ? (* src = "crypto_accelerator.v:237" *) _042_ : reg_6;
  assign _043_ = _020_ ? (* src = "crypto_accelerator.v:228" *) reg_14 : reg_4;
  assign _044_ = io_cyc ? (* src = "crypto_accelerator.v:227" *) _043_ : reg_4;
  assign _045_ = io_rev ? (* src = "crypto_accelerator.v:225" *) reg_6 : _044_;
  assign _010_ = io_enable ? (* src = "crypto_accelerator.v:224" *) _045_ : reg_5;
  assign _046_ = _019_ ? (* src = "crypto_accelerator.v:215" *) reg_14 : reg_3;
  assign _047_ = io_cyc ? (* src = "crypto_accelerator.v:214" *) _046_ : reg_3;
  assign _048_ = io_rev ? (* src = "crypto_accelerator.v:212" *) reg_5 : _047_;
  assign _009_ = io_enable ? (* src = "crypto_accelerator.v:211" *) _048_ : reg_4;
  assign _049_ = _018_ ? (* src = "crypto_accelerator.v:202" *) reg_14 : reg_2;
  assign _050_ = io_cyc ? (* src = "crypto_accelerator.v:201" *) _049_ : reg_2;
  assign _051_ = io_rev ? (* src = "crypto_accelerator.v:199" *) reg_4 : _050_;
  assign _008_ = io_enable ? (* src = "crypto_accelerator.v:198" *) _051_ : reg_3;
  assign _052_ = _017_ ? (* src = "crypto_accelerator.v:189" *) reg_14 : reg_1;
  assign _053_ = io_cyc ? (* src = "crypto_accelerator.v:188" *) _052_ : reg_1;
  assign _054_ = io_rev ? (* src = "crypto_accelerator.v:186" *) reg_3 : _053_;
  assign _007_ = io_enable ? (* src = "crypto_accelerator.v:185" *) _054_ : reg_2;
  assign _055_ = _016_ ? (* src = "crypto_accelerator.v:176" *) reg_14 : reg_0;
  assign _056_ = io_cyc ? (* src = "crypto_accelerator.v:175" *) _055_ : reg_0;
  assign _057_ = io_rev ? (* src = "crypto_accelerator.v:173" *) reg_2 : _056_;
  assign _006_ = io_enable ? (* src = "crypto_accelerator.v:172" *) _057_ : reg_1;
  assign _058_ = _015_ ? (* src = "crypto_accelerator.v:165" *) reg_14 : reg_0;
  assign _059_ = io_cyc ? (* src = "crypto_accelerator.v:164" *) _058_ : io_input;
  assign _060_ = io_rev ? (* src = "crypto_accelerator.v:162" *) reg_1 : _059_;
  assign _000_ = io_enable ? (* src = "crypto_accelerator.v:161" *) _060_ : reg_0;
  assign _T = io_tap ? (* src = "crypto_accelerator.v:71" *) 3'b000 : 3'b100;
  assign _GEN_75 = { 1'b0, _T };
  assign io_output_0 = reg_0;
  assign io_output_1 = reg_1;
  assign io_output_10 = reg_10;
  assign io_output_11 = reg_11;
  assign io_output_12 = reg_12;
  assign io_output_13 = reg_13;
  assign io_output_14 = reg_14;
  assign io_output_2 = reg_2;
  assign io_output_3 = reg_3;
  assign io_output_4 = reg_4;
  assign io_output_5 = reg_5;
  assign io_output_6 = reg_6;
  assign io_output_7 = reg_7;
  assign io_output_8 = reg_8;
  assign io_output_9 = reg_9;
endmodule
