module FP32_ADD_chn_a_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp32_add.v:363" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:364" *)
  output outsig;
  assign outsig = in_0;
endmodule
