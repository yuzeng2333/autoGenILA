module \$paramod\CDP_OCVT_mgc_in_wire_v1\rscid=5\width=2 (d, z);
  (* src = "./vmod/vlibs/HLS_cdp_ocvt.v:78" *)
  output [1:0] d;
  (* src = "./vmod/vlibs/HLS_cdp_ocvt.v:79" *)
  input [1:0] z;
  assign d = z;
endmodule
