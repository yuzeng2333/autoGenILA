module NV_NVDLA_RT_cmac_a2cacc(nvdla_core_clk, nvdla_core_rstn, mac2accu_src_pvld, mac2accu_src_mask, mac2accu_src_mode, mac2accu_src_data0, mac2accu_src_data1, mac2accu_src_data2, mac2accu_src_data3, mac2accu_src_data4, mac2accu_src_data5, mac2accu_src_data6, mac2accu_src_data7, mac2accu_src_pd, mac2accu_dst_pvld, mac2accu_dst_mask, mac2accu_dst_mode, mac2accu_dst_data0, mac2accu_dst_data1, mac2accu_dst_data2, mac2accu_dst_data3, mac2accu_dst_data4, mac2accu_dst_data5, mac2accu_dst_data6, mac2accu_dst_data7, mac2accu_dst_pd);
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:158" *)
  wire [131:0] _000_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:148" *)
  wire [43:0] _001_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:352" *)
  wire [131:0] _002_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:342" *)
  wire [43:0] _003_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:178" *)
  wire [131:0] _004_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:168" *)
  wire [43:0] _005_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:372" *)
  wire [131:0] _006_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:362" *)
  wire [43:0] _007_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:198" *)
  wire [131:0] _008_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:188" *)
  wire [43:0] _009_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:392" *)
  wire [131:0] _010_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:382" *)
  wire [43:0] _011_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:218" *)
  wire [131:0] _012_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:208" *)
  wire [43:0] _013_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:412" *)
  wire [131:0] _014_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:402" *)
  wire [43:0] _015_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:238" *)
  wire [131:0] _016_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:228" *)
  wire [43:0] _017_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:432" *)
  wire [131:0] _018_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:422" *)
  wire [43:0] _019_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:258" *)
  wire [131:0] _020_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:248" *)
  wire [43:0] _021_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:452" *)
  wire [131:0] _022_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:442" *)
  wire [43:0] _023_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:278" *)
  wire [131:0] _024_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:268" *)
  wire [43:0] _025_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:472" *)
  wire [131:0] _026_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:462" *)
  wire [43:0] _027_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:298" *)
  wire [131:0] _028_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:288" *)
  wire [43:0] _029_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:492" *)
  wire [131:0] _030_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:482" *)
  wire [43:0] _031_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:131" *)
  wire [7:0] _032_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:325" *)
  wire [7:0] _033_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:121" *)
  wire [8:0] _034_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:315" *)
  wire [8:0] _035_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:159" *)
  wire _036_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:179" *)
  wire _037_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:199" *)
  wire _038_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:219" *)
  wire _039_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:239" *)
  wire _040_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:259" *)
  wire _041_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:279" *)
  wire _042_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:299" *)
  wire _043_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:353" *)
  wire _044_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:373" *)
  wire _045_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:393" *)
  wire _046_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:413" *)
  wire _047_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:433" *)
  wire _048_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:453" *)
  wire _049_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:473" *)
  wire _050_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:493" *)
  wire _051_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:66" *)
  wire [175:0] mac2accu_data0_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:78" *)
  reg [175:0] mac2accu_data0_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:79" *)
  reg [175:0] mac2accu_data0_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:67" *)
  wire [175:0] mac2accu_data1_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:80" *)
  reg [175:0] mac2accu_data1_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:81" *)
  reg [175:0] mac2accu_data1_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:68" *)
  wire [175:0] mac2accu_data2_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:82" *)
  reg [175:0] mac2accu_data2_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:83" *)
  reg [175:0] mac2accu_data2_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:69" *)
  wire [175:0] mac2accu_data3_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:84" *)
  reg [175:0] mac2accu_data3_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:85" *)
  reg [175:0] mac2accu_data3_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:70" *)
  wire [175:0] mac2accu_data4_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:86" *)
  reg [175:0] mac2accu_data4_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:87" *)
  reg [175:0] mac2accu_data4_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:71" *)
  wire [175:0] mac2accu_data5_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:88" *)
  reg [175:0] mac2accu_data5_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:89" *)
  reg [175:0] mac2accu_data5_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:72" *)
  wire [175:0] mac2accu_data6_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:90" *)
  reg [175:0] mac2accu_data6_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:91" *)
  reg [175:0] mac2accu_data6_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:73" *)
  wire [175:0] mac2accu_data7_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:92" *)
  reg [175:0] mac2accu_data7_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:93" *)
  reg [175:0] mac2accu_data7_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:57" *)
  output [175:0] mac2accu_dst_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:58" *)
  output [175:0] mac2accu_dst_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:59" *)
  output [175:0] mac2accu_dst_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:60" *)
  output [175:0] mac2accu_dst_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:61" *)
  output [175:0] mac2accu_dst_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:62" *)
  output [175:0] mac2accu_dst_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:63" *)
  output [175:0] mac2accu_dst_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:64" *)
  output [175:0] mac2accu_dst_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:55" *)
  output [7:0] mac2accu_dst_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:56" *)
  output [7:0] mac2accu_dst_mode;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:65" *)
  output [8:0] mac2accu_dst_pd;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:54" *)
  output mac2accu_dst_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:74" *)
  wire [7:0] mac2accu_mask_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:94" *)
  reg [7:0] mac2accu_mask_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:95" *)
  reg [7:0] mac2accu_mask_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:75" *)
  wire [7:0] mac2accu_mode_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:96" *)
  reg [7:0] mac2accu_mode_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:97" *)
  reg [7:0] mac2accu_mode_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:76" *)
  wire [8:0] mac2accu_pd_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:98" *)
  reg [8:0] mac2accu_pd_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:99" *)
  reg [8:0] mac2accu_pd_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:77" *)
  wire mac2accu_pvld_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:100" *)
  reg mac2accu_pvld_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:101" *)
  reg mac2accu_pvld_d2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:45" *)
  input [175:0] mac2accu_src_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:46" *)
  input [175:0] mac2accu_src_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:47" *)
  input [175:0] mac2accu_src_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:48" *)
  input [175:0] mac2accu_src_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:49" *)
  input [175:0] mac2accu_src_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:50" *)
  input [175:0] mac2accu_src_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:51" *)
  input [175:0] mac2accu_src_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:52" *)
  input [175:0] mac2accu_src_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:43" *)
  input [7:0] mac2accu_src_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:44" *)
  input [7:0] mac2accu_src_mode;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:53" *)
  input [8:0] mac2accu_src_pd;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:42" *)
  input mac2accu_src_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:40" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:41" *)
  input nvdla_core_rstn;
  assign _036_ = mac2accu_src_mask[0] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:159" *) mac2accu_src_mode[0];
  assign _037_ = mac2accu_src_mask[1] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:179" *) mac2accu_src_mode[1];
  assign _038_ = mac2accu_src_mask[2] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:199" *) mac2accu_src_mode[2];
  assign _039_ = mac2accu_src_mask[3] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:219" *) mac2accu_src_mode[3];
  assign _040_ = mac2accu_src_mask[4] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:239" *) mac2accu_src_mode[4];
  assign _041_ = mac2accu_src_mask[5] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:259" *) mac2accu_src_mode[5];
  assign _042_ = mac2accu_src_mask[6] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:279" *) mac2accu_src_mode[6];
  assign _043_ = mac2accu_src_mask[7] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:299" *) mac2accu_src_mode[7];
  assign _044_ = mac2accu_mask_d1[0] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:353" *) mac2accu_mode_d1[0];
  assign _045_ = mac2accu_mask_d1[1] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:373" *) mac2accu_mode_d1[1];
  assign _046_ = mac2accu_mask_d1[2] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:393" *) mac2accu_mode_d1[2];
  assign _047_ = mac2accu_mask_d1[3] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:413" *) mac2accu_mode_d1[3];
  assign _048_ = mac2accu_mask_d1[4] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:433" *) mac2accu_mode_d1[4];
  assign _049_ = mac2accu_mask_d1[5] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:453" *) mac2accu_mode_d1[5];
  assign _050_ = mac2accu_mask_d1[6] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:473" *) mac2accu_mode_d1[6];
  assign _051_ = mac2accu_mask_d1[7] & (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:493" *) mac2accu_mode_d1[7];
  always @(posedge nvdla_core_clk)
      mac2accu_data7_d2[175:44] <= _030_;
  always @(posedge nvdla_core_clk)
      mac2accu_data7_d2[43:0] <= _031_;
  always @(posedge nvdla_core_clk)
      mac2accu_data6_d2[175:44] <= _026_;
  always @(posedge nvdla_core_clk)
      mac2accu_data6_d2[43:0] <= _027_;
  always @(posedge nvdla_core_clk)
      mac2accu_data5_d2[175:44] <= _022_;
  always @(posedge nvdla_core_clk)
      mac2accu_data5_d2[43:0] <= _023_;
  always @(posedge nvdla_core_clk)
      mac2accu_data4_d2[175:44] <= _018_;
  always @(posedge nvdla_core_clk)
      mac2accu_data4_d2[43:0] <= _019_;
  always @(posedge nvdla_core_clk)
      mac2accu_data3_d2[175:44] <= _014_;
  always @(posedge nvdla_core_clk)
      mac2accu_data3_d2[43:0] <= _015_;
  always @(posedge nvdla_core_clk)
      mac2accu_data2_d2[175:44] <= _010_;
  always @(posedge nvdla_core_clk)
      mac2accu_data2_d2[43:0] <= _011_;
  always @(posedge nvdla_core_clk)
      mac2accu_data1_d2[175:44] <= _006_;
  always @(posedge nvdla_core_clk)
      mac2accu_data1_d2[43:0] <= _007_;
  always @(posedge nvdla_core_clk)
      mac2accu_data0_d2[175:44] <= _002_;
  always @(posedge nvdla_core_clk)
      mac2accu_data0_d2[43:0] <= _003_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mac2accu_mask_d2 <= 8'b00000000;
    else
      mac2accu_mask_d2 <= mac2accu_mask_d1;
  always @(posedge nvdla_core_clk)
      mac2accu_mode_d2 <= _033_;
  always @(posedge nvdla_core_clk)
      mac2accu_pd_d2 <= _035_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mac2accu_pvld_d2 <= 1'b0;
    else
      mac2accu_pvld_d2 <= mac2accu_pvld_d1;
  always @(posedge nvdla_core_clk)
      mac2accu_data7_d1[175:44] <= _028_;
  always @(posedge nvdla_core_clk)
      mac2accu_data7_d1[43:0] <= _029_;
  always @(posedge nvdla_core_clk)
      mac2accu_data6_d1[175:44] <= _024_;
  always @(posedge nvdla_core_clk)
      mac2accu_data6_d1[43:0] <= _025_;
  always @(posedge nvdla_core_clk)
      mac2accu_data5_d1[175:44] <= _020_;
  always @(posedge nvdla_core_clk)
      mac2accu_data5_d1[43:0] <= _021_;
  always @(posedge nvdla_core_clk)
      mac2accu_data4_d1[175:44] <= _016_;
  always @(posedge nvdla_core_clk)
      mac2accu_data4_d1[43:0] <= _017_;
  always @(posedge nvdla_core_clk)
      mac2accu_data3_d1[175:44] <= _012_;
  always @(posedge nvdla_core_clk)
      mac2accu_data3_d1[43:0] <= _013_;
  always @(posedge nvdla_core_clk)
      mac2accu_data2_d1[175:44] <= _008_;
  always @(posedge nvdla_core_clk)
      mac2accu_data2_d1[43:0] <= _009_;
  always @(posedge nvdla_core_clk)
      mac2accu_data1_d1[175:44] <= _004_;
  always @(posedge nvdla_core_clk)
      mac2accu_data1_d1[43:0] <= _005_;
  always @(posedge nvdla_core_clk)
      mac2accu_data0_d1[175:44] <= _000_;
  always @(posedge nvdla_core_clk)
      mac2accu_data0_d1[43:0] <= _001_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mac2accu_mask_d1 <= 8'b00000000;
    else
      mac2accu_mask_d1 <= mac2accu_src_mask;
  always @(posedge nvdla_core_clk)
      mac2accu_mode_d1 <= _032_;
  always @(posedge nvdla_core_clk)
      mac2accu_pd_d1 <= _034_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mac2accu_pvld_d1 <= 1'b0;
    else
      mac2accu_pvld_d1 <= mac2accu_src_pvld;
  assign _030_ = _051_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:493" *) mac2accu_data7_d1[175:44] : mac2accu_data7_d2[175:44];
  assign _031_ = mac2accu_mask_d1[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:483" *) mac2accu_data7_d1[43:0] : mac2accu_data7_d2[43:0];
  assign _026_ = _050_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:473" *) mac2accu_data6_d1[175:44] : mac2accu_data6_d2[175:44];
  assign _027_ = mac2accu_mask_d1[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:463" *) mac2accu_data6_d1[43:0] : mac2accu_data6_d2[43:0];
  assign _022_ = _049_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:453" *) mac2accu_data5_d1[175:44] : mac2accu_data5_d2[175:44];
  assign _023_ = mac2accu_mask_d1[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:443" *) mac2accu_data5_d1[43:0] : mac2accu_data5_d2[43:0];
  assign _018_ = _048_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:433" *) mac2accu_data4_d1[175:44] : mac2accu_data4_d2[175:44];
  assign _019_ = mac2accu_mask_d1[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:423" *) mac2accu_data4_d1[43:0] : mac2accu_data4_d2[43:0];
  assign _014_ = _047_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:413" *) mac2accu_data3_d1[175:44] : mac2accu_data3_d2[175:44];
  assign _015_ = mac2accu_mask_d1[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:403" *) mac2accu_data3_d1[43:0] : mac2accu_data3_d2[43:0];
  assign _010_ = _046_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:393" *) mac2accu_data2_d1[175:44] : mac2accu_data2_d2[175:44];
  assign _011_ = mac2accu_mask_d1[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:383" *) mac2accu_data2_d1[43:0] : mac2accu_data2_d2[43:0];
  assign _006_ = _045_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:373" *) mac2accu_data1_d1[175:44] : mac2accu_data1_d2[175:44];
  assign _007_ = mac2accu_mask_d1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:363" *) mac2accu_data1_d1[43:0] : mac2accu_data1_d2[43:0];
  assign _002_ = _044_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:353" *) mac2accu_data0_d1[175:44] : mac2accu_data0_d2[175:44];
  assign _003_ = mac2accu_mask_d1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:343" *) mac2accu_data0_d1[43:0] : mac2accu_data0_d2[43:0];
  assign _033_ = mac2accu_pvld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:326" *) mac2accu_mode_d1 : mac2accu_mode_d2;
  assign _035_ = mac2accu_pvld_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:316" *) mac2accu_pd_d1 : mac2accu_pd_d2;
  assign _028_ = _043_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:299" *) mac2accu_src_data7[175:44] : mac2accu_data7_d1[175:44];
  assign _029_ = mac2accu_src_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:289" *) mac2accu_src_data7[43:0] : mac2accu_data7_d1[43:0];
  assign _024_ = _042_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:279" *) mac2accu_src_data6[175:44] : mac2accu_data6_d1[175:44];
  assign _025_ = mac2accu_src_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:269" *) mac2accu_src_data6[43:0] : mac2accu_data6_d1[43:0];
  assign _020_ = _041_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:259" *) mac2accu_src_data5[175:44] : mac2accu_data5_d1[175:44];
  assign _021_ = mac2accu_src_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:249" *) mac2accu_src_data5[43:0] : mac2accu_data5_d1[43:0];
  assign _016_ = _040_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:239" *) mac2accu_src_data4[175:44] : mac2accu_data4_d1[175:44];
  assign _017_ = mac2accu_src_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:229" *) mac2accu_src_data4[43:0] : mac2accu_data4_d1[43:0];
  assign _012_ = _039_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:219" *) mac2accu_src_data3[175:44] : mac2accu_data3_d1[175:44];
  assign _013_ = mac2accu_src_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:209" *) mac2accu_src_data3[43:0] : mac2accu_data3_d1[43:0];
  assign _008_ = _038_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:199" *) mac2accu_src_data2[175:44] : mac2accu_data2_d1[175:44];
  assign _009_ = mac2accu_src_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:189" *) mac2accu_src_data2[43:0] : mac2accu_data2_d1[43:0];
  assign _004_ = _037_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:179" *) mac2accu_src_data1[175:44] : mac2accu_data1_d1[175:44];
  assign _005_ = mac2accu_src_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:169" *) mac2accu_src_data1[43:0] : mac2accu_data1_d1[43:0];
  assign _000_ = _036_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:159" *) mac2accu_src_data0[175:44] : mac2accu_data0_d1[175:44];
  assign _001_ = mac2accu_src_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:149" *) mac2accu_src_data0[43:0] : mac2accu_data0_d1[43:0];
  assign _032_ = mac2accu_src_pvld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:132" *) mac2accu_src_mode : mac2accu_mode_d1;
  assign _034_ = mac2accu_src_pvld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_cmac_a2cacc.v:122" *) mac2accu_src_pd : mac2accu_pd_d1;
  assign mac2accu_data0_d0 = mac2accu_src_data0;
  assign mac2accu_data1_d0 = mac2accu_src_data1;
  assign mac2accu_data2_d0 = mac2accu_src_data2;
  assign mac2accu_data3_d0 = mac2accu_src_data3;
  assign mac2accu_data4_d0 = mac2accu_src_data4;
  assign mac2accu_data5_d0 = mac2accu_src_data5;
  assign mac2accu_data6_d0 = mac2accu_src_data6;
  assign mac2accu_data7_d0 = mac2accu_src_data7;
  assign mac2accu_dst_data0 = mac2accu_data0_d2;
  assign mac2accu_dst_data1 = mac2accu_data1_d2;
  assign mac2accu_dst_data2 = mac2accu_data2_d2;
  assign mac2accu_dst_data3 = mac2accu_data3_d2;
  assign mac2accu_dst_data4 = mac2accu_data4_d2;
  assign mac2accu_dst_data5 = mac2accu_data5_d2;
  assign mac2accu_dst_data6 = mac2accu_data6_d2;
  assign mac2accu_dst_data7 = mac2accu_data7_d2;
  assign mac2accu_dst_mask = mac2accu_mask_d2;
  assign mac2accu_dst_mode = mac2accu_mode_d2;
  assign mac2accu_dst_pd = mac2accu_pd_d2;
  assign mac2accu_dst_pvld = mac2accu_pvld_d2;
  assign mac2accu_mask_d0 = mac2accu_src_mask;
  assign mac2accu_mode_d0 = mac2accu_src_mode;
  assign mac2accu_pd_d0 = mac2accu_src_pd;
  assign mac2accu_pvld_d0 = mac2accu_src_pvld;
endmodule
