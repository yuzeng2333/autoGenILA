module \$paramod\SDP_X_mgc_in_wire_v1\rscid=19\width=1 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:109" *)
  output d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:110" *)
  input z;
  assign d = z;
endmodule
