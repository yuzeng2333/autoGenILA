module FP32_SUB_chn_a_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp32_sub.v:363" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp32_sub.v:364" *)
  output outsig;
  assign outsig = in_0;
endmodule
