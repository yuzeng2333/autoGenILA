module \$paramod\CDMA_mgc_in_wire_v1\rscid=3\width=16 (d, z);
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:78" *)
  output [15:0] d;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_CVT_cell.v:79" *)
  input [15:0] z;
  assign d = z;
endmodule
