module NV_NVDLA_SDP_CORE_Y_idx_core(nvdla_core_clk, nvdla_core_rstn, chn_lut_in_rsc_z, chn_lut_in_rsc_vz, chn_lut_in_rsc_lz, cfg_lut_le_start_rsc_z, cfg_lut_lo_start_rsc_z, cfg_lut_le_index_offset_rsc_z, cfg_lut_le_index_select_rsc_z, cfg_lut_lo_index_select_rsc_z, cfg_lut_le_function_rsc_z, cfg_lut_uflow_priority_rsc_z, cfg_lut_oflow_priority_rsc_z, cfg_lut_hybrid_priority_rsc_z, cfg_precision_rsc_z, chn_lut_out_rsc_z, chn_lut_out_rsc_vz, chn_lut_out_rsc_lz, chn_lut_in_rsci_oswt, chn_lut_in_rsci_oswt_unreg, chn_lut_out_rsci_oswt, chn_lut_out_rsci_oswt_unreg);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13452" *)
  wire _00039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13605" *)
  wire [7:0] _00040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13605" *)
  wire [7:0] _00041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13605" *)
  wire [7:0] _00042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13605" *)
  wire [7:0] _00043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13605" *)
  wire [7:0] _00044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13605" *)
  wire [7:0] _00045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13622" *)
  wire [8:0] _00061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13771" *)
  wire [8:0] _00062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13771" *)
  wire [8:0] _00063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13771" *)
  wire [8:0] _00064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13771" *)
  wire [8:0] _00065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13777" *)
  wire [7:0] _00066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13777" *)
  wire [7:0] _00067_;
  wire [22:0] _00068_;
  wire [22:0] _00069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13723" *)
  wire [34:0] _00089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10082" *)
  wire [7:0] _00090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire [7:0] _00091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire [7:0] _00092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire [7:0] _00093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8282" *)
  wire [49:0] _00094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8337" *)
  wire [49:0] _00095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8378" *)
  wire [49:0] _00096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8427" *)
  wire [49:0] _00097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10122" *)
  wire _00098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10122" *)
  wire _00099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10122" *)
  wire _00100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10122" *)
  wire _00101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8641" *)
  wire _00102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8794" *)
  wire _00103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8794" *)
  wire _00104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8794" *)
  wire _00105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10303" *)
  wire _00106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8564" *)
  wire _00107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11407" *)
  wire _00108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11371" *)
  wire _00109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10325" *)
  wire _00110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8784" *)
  wire _00111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11425" *)
  wire _00112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10347" *)
  wire _00113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8933" *)
  wire _00114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11453" *)
  wire _00115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10369" *)
  wire _00116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9053" *)
  wire _00117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10082" *)
  wire [7:0] _00118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire [7:0] _00119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire [7:0] _00120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire [7:0] _00121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8144" *)
  wire [7:0] _00122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10093" *)
  wire [7:0] _00123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10208" *)
  wire [7:0] _00124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10226" *)
  wire [7:0] _00125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8306" *)
  wire [49:0] _00126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8359" *)
  wire [49:0] _00127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8408" *)
  wire [49:0] _00128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8439" *)
  wire [49:0] _00129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10155" *)
  wire _00130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10155" *)
  wire _00131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10155" *)
  wire _00132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10155" *)
  wire _00133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8701" *)
  wire _00134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8701" *)
  wire _00135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8701" *)
  wire _00136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8701" *)
  wire _00137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10314" *)
  wire _00138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8691" *)
  wire _00139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11416" *)
  wire _00140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11398" *)
  wire _00141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10336" *)
  wire _00142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8857" *)
  wire _00143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11434" *)
  wire _00144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10358" *)
  wire _00145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8977" *)
  wire _00146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11480" *)
  wire _00147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10380" *)
  wire _00148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9097" *)
  wire _00149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8671" *)
  wire [7:0] _00150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8830" *)
  wire [7:0] _00151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8964" *)
  wire [7:0] _00152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9084" *)
  wire [7:0] _00153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10785" *)
  wire [22:0] _00154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10917" *)
  wire [22:0] _00155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11025" *)
  wire [22:0] _00156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11151" *)
  wire [22:0] _00157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8144" *)
  wire [7:0] _00158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8294" *)
  wire [7:0] _00159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10093" *)
  wire [7:0] _00160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8349" *)
  wire [7:0] _00161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10104" *)
  wire [7:0] _00162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8390" *)
  wire [7:0] _00163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10113" *)
  wire [7:0] _00164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8390" *)
  wire [7:0] _00165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9289" *)
  wire _00166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9349" *)
  wire _00167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9409" *)
  wire _00168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9229" *)
  wire _00169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9683" *)
  wire [255:0] _00170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9801" *)
  wire [255:0] _00171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9889" *)
  wire [255:0] _00172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9977" *)
  wire [255:0] _00173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9269" *)
  wire _00174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9329" *)
  wire _00175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9389" *)
  wire _00176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9209" *)
  wire _00177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9621" *)
  wire [255:0] _00178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9751" *)
  wire [255:0] _00179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9845" *)
  wire [255:0] _00180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9943" *)
  wire [255:0] _00181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8531" *)
  wire _00182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8751" *)
  wire _00183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8899" *)
  wire _00184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9019" *)
  wire _00185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8660" *)
  wire _00186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8819" *)
  wire _00187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8953" *)
  wire _00188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9073" *)
  wire _00189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11223" *)
  wire [30:0] _00190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11247" *)
  wire [30:0] _00191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11275" *)
  wire [30:0] _00192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11291" *)
  wire [30:0] _00193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10616" *)
  wire _00194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9675" *)
  wire _00195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10596" *)
  wire _00196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9793" *)
  wire _00197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10568" *)
  wire _00198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9881" *)
  wire _00199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10548" *)
  wire _00200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9969" *)
  wire _00201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10140" *)
  wire _00202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10249" *)
  wire _00203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8499" *)
  wire _00204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10264" *)
  wire _00206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8719" *)
  wire _00207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10264" *)
  wire _00208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8867" *)
  wire _00209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10249" *)
  wire _00211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8987" *)
  wire _00212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11470" *)
  wire _00222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11388" *)
  wire _00223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10278" *)
  wire _00224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10234" *)
  wire _00225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10234" *)
  wire _00226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10234" *)
  wire _00227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11462" *)
  wire _00228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11380" *)
  wire _00229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10511" *)
  wire _00230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9613" *)
  wire _00231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10499" *)
  wire _00232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9743" *)
  wire _00233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10487" *)
  wire _00234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9837" *)
  wire _00235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10455" *)
  wire _00236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9935" *)
  wire _00237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10249" *)
  wire _00238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8144" *)
  wire _00240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8294" *)
  wire _00241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10288" *)
  wire _00243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8843" *)
  wire _00244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8349" *)
  wire _00245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8843" *)
  wire _00246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10288" *)
  wire _00247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8390" *)
  wire _00250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10288" *)
  wire _00252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11443" *)
  wire _00255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11489" *)
  wire _00256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8294" *)
  wire _00257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8843" *)
  wire _00259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8390" *)
  wire _00260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8390" *)
  wire _00262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11443" *)
  wire _00264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11489" *)
  wire _00265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire _00267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire _00268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire _00270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire _00273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire [7:0] _00274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire [7:0] _00275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire [7:0] _00276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9115" *)
  wire [7:0] _00277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire [7:0] _00278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire [7:0] _00279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire [7:0] _00280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire [30:0] _00281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire [30:0] _00282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire [31:0] _00283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire [7:0] _00284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire [7:0] _00285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire [7:0] _00286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire [30:0] _00287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8683" *)
  wire [30:0] _00288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire [31:0] _00289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire _00291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire _00292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire _00294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire _00296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire _00297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire _00299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10695" *)
  wire [1:0] _00300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [1:0] _00301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire [1:0] _00302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [1:0] _00303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9649" *)
  wire [1:0] _00304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7880" *)
  wire _00305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7890" *)
  wire _00306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [22:0] _00307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [11:0] _00308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [11:0] _00309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [22:0] _00310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [127:0] _00311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7998" *)
  wire _00316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8019" *)
  wire _00317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8040" *)
  wire _00318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8061" *)
  wire _00319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7998" *)
  wire _00320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8019" *)
  wire _00321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8040" *)
  wire _00322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8061" *)
  wire _00323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [5:0] _00324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7998" *)
  wire _00325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7998" *)
  wire _00326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7998" *)
  wire _00327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [5:0] _00328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8019" *)
  wire _00329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8019" *)
  wire _00330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8019" *)
  wire _00331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [5:0] _00332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8040" *)
  wire _00333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8040" *)
  wire _00334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8040" *)
  wire _00335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [5:0] _00336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8061" *)
  wire _00337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8061" *)
  wire _00338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8061" *)
  wire _00339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire _00347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [22:0] _00348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [11:0] _00349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [22:0] _00350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [11:0] _00351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7880" *)
  wire _00352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire [127:0] _00353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire [127:0] _00354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire [127:0] _00355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [127:0] _00356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [127:0] _00357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10140" *)
  wire _00358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10140" *)
  wire _00359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8144" *)
  wire _00360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9229" *)
  wire [7:0] _00361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9665" *)
  wire _00362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9209" *)
  wire [7:0] _00363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9603" *)
  wire _00364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8531" *)
  wire [22:0] _00365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8650" *)
  wire [22:0] _00367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10685" *)
  wire [1:0] _00368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10795" *)
  wire [31:0] _00370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11333" *)
  wire _00371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10578" *)
  wire _00372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9239" *)
  wire _00373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10823" *)
  wire _00374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10703" *)
  wire [31:0] _00375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9123" *)
  wire _00376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11499" *)
  wire [5:0] _00377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire _00378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire _00379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10654" *)
  wire _00381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9143" *)
  wire _00382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9289" *)
  wire [7:0] _00386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9783" *)
  wire _00387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9269" *)
  wire [7:0] _00388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9733" *)
  wire _00389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8751" *)
  wire [22:0] _00390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8843" *)
  wire _00391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8809" *)
  wire [22:0] _00392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10869" *)
  wire [1:0] _00393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10927" *)
  wire [31:0] _00395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11333" *)
  wire _00396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10578" *)
  wire _00397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9299" *)
  wire _00398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10955" *)
  wire _00399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10879" *)
  wire [31:0] _00400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9249" *)
  wire _00401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11527" *)
  wire [5:0] _00402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire _00403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire _00404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10654" *)
  wire _00406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9143" *)
  wire _00407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10200" *)
  wire _00410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9349" *)
  wire [7:0] _00411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9871" *)
  wire _00412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9329" *)
  wire [7:0] _00413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9827" *)
  wire _00414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8899" *)
  wire [22:0] _00415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8943" *)
  wire [22:0] _00417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10989" *)
  wire [1:0] _00418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11035" *)
  wire [31:0] _00420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11333" *)
  wire _00421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10530" *)
  wire _00422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9359" *)
  wire _00423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11063" *)
  wire _00424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10999" *)
  wire [31:0] _00425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9309" *)
  wire _00426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11555" *)
  wire [5:0] _00427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire _00428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire _00429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10654" *)
  wire _00431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9143" *)
  wire _00432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10216" *)
  wire _00435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10216" *)
  wire _00436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9409" *)
  wire [7:0] _00437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9959" *)
  wire _00438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9389" *)
  wire [7:0] _00439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9925" *)
  wire _00440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9019" *)
  wire [22:0] _00441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9063" *)
  wire [22:0] _00443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11115" *)
  wire [1:0] _00444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11161" *)
  wire [31:0] _00446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11333" *)
  wire _00447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10530" *)
  wire _00448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9419" *)
  wire _00449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11189" *)
  wire _00450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11125" *)
  wire [31:0] _00451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9369" *)
  wire _00452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11583" *)
  wire [5:0] _00453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire _00454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire _00455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11107" *)
  wire _00457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9143" *)
  wire _00458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10399" *)
  wire [31:0] _00459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11519" *)
  wire [31:0] _00460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10415" *)
  wire [31:0] _00461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11547" *)
  wire [31:0] _00462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10431" *)
  wire [31:0] _00463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11575" *)
  wire [31:0] _00464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10447" *)
  wire [31:0] _00465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11603" *)
  wire [31:0] _00466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10003" *)
  wire _00467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10037" *)
  wire _00468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10037" *)
  wire _00469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10003" *)
  wire _00470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11681" *)
  wire _00471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11619" *)
  wire _00472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11325" *)
  wire _00473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10833" *)
  wire _00474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11669" *)
  wire _00475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11635" *)
  wire _00476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11315" *)
  wire _00477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10965" *)
  wire _00478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11669" *)
  wire _00479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11635" *)
  wire _00480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11315" *)
  wire _00481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11073" *)
  wire _00482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11669" *)
  wire _00483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11661" *)
  wire _00484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11307" *)
  wire _00485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11073" *)
  wire _00486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9715" *)
  wire _00487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9809" *)
  wire _00488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9907" *)
  wire _00489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9585" *)
  wire _00490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11239" *)
  wire _00491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10769" *)
  wire _00492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9219" *)
  wire _00493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11267" *)
  wire _00494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10897" *)
  wire _00495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9279" *)
  wire _00496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11283" *)
  wire _00497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11017" *)
  wire _00498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9339" *)
  wire _00499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11299" *)
  wire _00500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11143" *)
  wire _00501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9399" *)
  wire _00502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10391" *)
  wire [31:0] _00503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11511" *)
  wire [31:0] _00504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10407" *)
  wire [31:0] _00505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11539" *)
  wire [31:0] _00506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10423" *)
  wire [31:0] _00507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11567" *)
  wire [31:0] _00508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10439" *)
  wire [31:0] _00509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11595" *)
  wire [31:0] _00510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10019" *)
  wire _00511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10053" *)
  wire _00512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10019" *)
  wire _00513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10019" *)
  wire _00514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11231" *)
  wire _00515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10777" *)
  wire _00516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11255" *)
  wire _00517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10905" *)
  wire _00518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11255" *)
  wire _00519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10905" *)
  wire _00520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11255" *)
  wire _00521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10905" *)
  wire _00522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9595" *)
  wire [34:0] _00523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9725" *)
  wire [34:0] _00524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9819" *)
  wire [34:0] _00525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9917" *)
  wire [34:0] _00526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10467" *)
  wire _00527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9853" *)
  wire _00528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9637" *)
  wire _00529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10522" *)
  wire _00530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9629" *)
  wire _00531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9637" *)
  wire _00532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10467" *)
  wire _00533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9759" *)
  wire _00534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9767" *)
  wire _00535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10467" *)
  wire _00536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9853" *)
  wire _00537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9637" *)
  wire _00538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11199" *)
  wire _00539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11199" *)
  wire _00540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11199" *)
  wire _00541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11214" *)
  wire _00542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10479" *)
  wire _00543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire _00545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9657" *)
  wire [34:0] _00546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9775" *)
  wire [34:0] _00547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9863" *)
  wire [34:0] _00548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9951" *)
  wire [34:0] _00549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10558" *)
  wire _00550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9897" *)
  wire _00551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9701" *)
  wire _00552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10606" *)
  wire _00553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9691" *)
  wire _00554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9701" *)
  wire _00555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10606" *)
  wire _00556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9691" *)
  wire _00557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9701" *)
  wire _00558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10558" *)
  wire _00559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9897" *)
  wire _00560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9701" *)
  wire _00561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10638" *)
  wire _00562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10841" *)
  wire _00563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10973" *)
  wire _00564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11091" *)
  wire _00565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11611" *)
  wire [30:0] _00566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11627" *)
  wire [30:0] _00567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11645" *)
  wire [30:0] _00568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11653" *)
  wire [30:0] _00569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10646" *)
  wire _00571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9135" *)
  wire _00572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10849" *)
  wire _00574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9261" *)
  wire _00575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10981" *)
  wire _00577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9321" *)
  wire _00578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8457" *)
  wire _00579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11099" *)
  wire _00580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9381" *)
  wire _00581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11083" *)
  wire _00582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10626" *)
  wire _00583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10626" *)
  wire _00584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10626" *)
  wire _00585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [22:0] _00586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [22:0] _00589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [22:0] _00592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [22:0] _00595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [5:0] _00617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9985" *)
  wire _00618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9985" *)
  wire _00619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9985" *)
  wire _00620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9985" *)
  wire _00621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire [34:0] _00625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11333" *)
  wire [7:0] _00626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10578" *)
  wire [7:0] _00627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10037" *)
  wire [7:0] _00628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11333" *)
  wire [7:0] _00629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10578" *)
  wire [7:0] _00630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10037" *)
  wire [7:0] _00631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11333" *)
  wire [7:0] _00632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10530" *)
  wire [7:0] _00633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10003" *)
  wire [7:0] _00634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11333" *)
  wire [7:0] _00635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10530" *)
  wire [7:0] _00636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10003" *)
  wire [7:0] _00637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10064" *)
  wire _00638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10064" *)
  wire _00640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10064" *)
  wire _00642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10064" *)
  wire _00644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8090" *)
  wire _00647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8220" *)
  wire _00648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8449" *)
  wire _00649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9107" *)
  wire _00650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9429" *)
  wire _00651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8554" *)
  wire [5:0] _00652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8543" *)
  wire [1:0] _00653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8774" *)
  wire [5:0] _00654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8763" *)
  wire [1:0] _00655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8923" *)
  wire [5:0] _00656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8911" *)
  wire [1:0] _00657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9043" *)
  wire [5:0] _00658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9031" *)
  wire [1:0] _00659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8273" *)
  wire [5:0] _00660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8264" *)
  wire [1:0] _00661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8328" *)
  wire [5:0] _00662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8316" *)
  wire [1:0] _00663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8369" *)
  wire [5:0] _00664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8316" *)
  wire [1:0] _00665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8418" *)
  wire [5:0] _00666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8316" *)
  wire [1:0] _00667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10677" *)
  wire [22:0] _00668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10666" *)
  wire [7:0] _00669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10749" *)
  wire [22:0] _00670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10857" *)
  wire [7:0] _00671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10749" *)
  wire [22:0] _00672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10749" *)
  wire [22:0] _00673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10857" *)
  wire [7:0] _00674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10857" *)
  wire [7:0] _00675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8390" *)
  wire _00677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire _00678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire _00679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8098" *)
  wire [1:0] _00680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8228" *)
  wire [1:0] _00681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8082" *)
  wire _00682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8134" *)
  wire _00683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8144" *)
  wire _00684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10814" *)
  wire [7:0] _00686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10804" *)
  wire _00687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10726" *)
  wire _00688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10740" *)
  wire [2:0] _00689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10749" *)
  wire [3:0] _00690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10712" *)
  wire _00691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8520" *)
  wire [1:0] _00692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8510" *)
  wire _00693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10946" *)
  wire [7:0] _00697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10936" *)
  wire _00698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10726" *)
  wire _00699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10888" *)
  wire [2:0] _00700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10749" *)
  wire [3:0] _00701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10712" *)
  wire _00702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8740" *)
  wire [1:0] _00703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8730" *)
  wire _00704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11054" *)
  wire [7:0] _00708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11044" *)
  wire _00709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10726" *)
  wire _00710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11008" *)
  wire [2:0] _00711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10749" *)
  wire [3:0] _00712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10712" *)
  wire _00713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8888" *)
  wire [1:0] _00714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8878" *)
  wire _00715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire _00717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8603" *)
  wire _00718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11180" *)
  wire [7:0] _00719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11170" *)
  wire _00720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10726" *)
  wire _00721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11134" *)
  wire [2:0] _00722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10749" *)
  wire [3:0] _00723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10712" *)
  wire _00724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9008" *)
  wire [1:0] _00725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8998" *)
  wire _00726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9437" *)
  wire _00727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10064" *)
  wire _00728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10064" *)
  wire _00729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10064" *)
  wire _00730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10064" *)
  wire _00731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10122" *)
  wire _00732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10122" *)
  wire _00733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10122" *)
  wire _00734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10122" *)
  wire _00735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10140" *)
  wire _00736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10140" *)
  wire _00737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10140" *)
  wire _00738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10155" *)
  wire _00739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10155" *)
  wire _00740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10155" *)
  wire _00741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10155" *)
  wire _00742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10173" *)
  wire _00749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10234" *)
  wire _00750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10234" *)
  wire _00751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10234" *)
  wire _00752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10249" *)
  wire _00753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10249" *)
  wire _00754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10249" *)
  wire _00755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10278" *)
  wire _00756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10288" *)
  wire _00757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10288" *)
  wire _00758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10288" *)
  wire _00759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10548" *)
  wire _00760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10568" *)
  wire _00761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10596" *)
  wire _00762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10616" *)
  wire _00763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11199" *)
  wire _00764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11199" *)
  wire _00765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11199" *)
  wire _00766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11214" *)
  wire _00767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11371" *)
  wire _00768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11388" *)
  wire _00769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11398" *)
  wire _00770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11407" *)
  wire _00771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11416" *)
  wire _00772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11425" *)
  wire _00773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11434" *)
  wire _00774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11453" *)
  wire _00775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11470" *)
  wire _00776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11480" *)
  wire _00777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7998" *)
  wire _00778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7998" *)
  wire _00779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7998" *)
  wire _00780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7998" *)
  wire _00781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7998" *)
  wire _00782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8019" *)
  wire _00783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8019" *)
  wire _00784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8019" *)
  wire _00785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8019" *)
  wire _00786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8019" *)
  wire _00787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8040" *)
  wire _00788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8040" *)
  wire _00789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8040" *)
  wire _00790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8040" *)
  wire _00791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8040" *)
  wire _00792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8061" *)
  wire _00793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8061" *)
  wire _00794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8061" *)
  wire _00795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8061" *)
  wire _00796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8061" *)
  wire _00797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8564" *)
  wire _00798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8573" *)
  wire _00806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8641" *)
  wire _00807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8660" *)
  wire _00808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8691" *)
  wire _00809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8701" *)
  wire _00810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8701" *)
  wire _00811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8701" *)
  wire _00812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8701" *)
  wire _00813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8784" *)
  wire _00814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8794" *)
  wire _00815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8794" *)
  wire _00816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8794" *)
  wire _00817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8819" *)
  wire _00818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8857" *)
  wire _00819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8933" *)
  wire _00820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8953" *)
  wire _00821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8977" *)
  wire _00822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9053" *)
  wire _00823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9073" *)
  wire _00824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9097" *)
  wire _00825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9123" *)
  wire _00826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9219" *)
  wire _00827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9249" *)
  wire _00828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9279" *)
  wire _00829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9309" *)
  wire _00830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9339" *)
  wire _00831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9369" *)
  wire _00832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9399" *)
  wire _00833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9585" *)
  wire _00834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9715" *)
  wire _00835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9809" *)
  wire _00836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9907" *)
  wire _00837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9985" *)
  wire _00838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9985" *)
  wire _00839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9985" *)
  wire _00840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9985" *)
  wire _00841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [11:0] _00842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [11:0] _00843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [11:0] _00844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7898" *)
  wire [11:0] _00845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10785" *)
  wire [22:0] _00846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10917" *)
  wire [22:0] _00847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11025" *)
  wire [22:0] _00848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11151" *)
  wire [22:0] _00849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8306" *)
  wire [49:0] _00850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8359" *)
  wire [49:0] _00851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8408" *)
  wire [49:0] _00852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8439" *)
  wire [49:0] _00853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11499" *)
  wire [5:0] _00854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11527" *)
  wire [5:0] _00855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11555" *)
  wire [5:0] _00856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11583" *)
  wire [5:0] _00857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9157" *)
  wire [5:0] _00861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10082" *)
  wire [7:0] _00862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10093" *)
  wire [7:0] _00863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10104" *)
  wire [7:0] _00864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10113" *)
  wire [7:0] _00865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8144" *)
  wire [7:0] _00866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire [7:0] _00867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire [7:0] _00868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8163" *)
  wire [7:0] _00869_;
  wire [49:0] _00870_;
  wire [49:0] _00871_;
  wire [49:0] _00872_;
  wire [49:0] _00873_;
  wire [49:0] _00874_;
  wire [49:0] _00875_;
  wire [49:0] _00876_;
  wire [49:0] _00877_;
  wire [49:0] _00878_;
  wire [49:0] _00879_;
  wire [49:0] _00880_;
  wire [49:0] _00881_;
  wire [7:0] _00882_;
  wire [7:0] _00883_;
  wire [7:0] _00884_;
  wire [7:0] _00885_;
  wire [7:0] _00886_;
  wire [7:0] _00887_;
  wire [7:0] _00888_;
  wire [7:0] _00889_;
  wire [8:0] _00890_;
  wire [8:0] _00891_;
  wire [8:0] _00892_;
  wire [8:0] _00893_;
  wire [8:0] _00894_;
  wire [8:0] _00895_;
  wire [8:0] _00896_;
  wire [8:0] _00897_;
  wire [23:0] _00898_;
  wire [23:0] _00899_;
  wire [23:0] _00900_;
  wire [23:0] _00901_;
  wire [8:0] _00902_;
  wire [8:0] _00903_;
  wire [8:0] _00904_;
  wire [8:0] _00905_;
  wire [8:0] _00906_;
  wire [8:0] _00907_;
  wire [8:0] _00908_;
  wire [8:0] _00909_;
  wire [23:0] _00910_;
  wire [23:0] _00911_;
  wire [23:0] _00912_;
  wire [23:0] _00913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10013" *)
  wire _00914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10016" *)
  wire _00915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10047" *)
  wire _00916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10050" *)
  wire _00917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10057" *)
  wire _00918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10058" *)
  wire _00919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10108" *)
  wire _00920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10108" *)
  wire _00921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10117" *)
  wire _00922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10117" *)
  wire _00923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10204" *)
  wire _00924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10204" *)
  wire _00925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10212" *)
  wire _00926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10230" *)
  wire _00927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10282" *)
  wire _00928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10283" *)
  wire _00929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10308" *)
  wire _00930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10308" *)
  wire _00931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10319" *)
  wire _00932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10319" *)
  wire _00933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10330" *)
  wire _00934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10330" *)
  wire _00935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10341" *)
  wire _00936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10341" *)
  wire _00937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10352" *)
  wire _00938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10352" *)
  wire _00939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10363" *)
  wire _00940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10363" *)
  wire _00941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10374" *)
  wire _00942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10374" *)
  wire _00943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10385" *)
  wire _00944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10385" *)
  wire _00945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10395" *)
  wire _00946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10403" *)
  wire _00947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10411" *)
  wire _00948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10419" *)
  wire _00949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10427" *)
  wire _00950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10435" *)
  wire _00951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10443" *)
  wire _00952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10451" *)
  wire _00953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10459" *)
  wire _00954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10460" *)
  wire _00955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10483" *)
  wire _00956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10492" *)
  wire _00957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10504" *)
  wire _00958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10516" *)
  wire _00959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10526" *)
  wire _00960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10552" *)
  wire _00961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10553" *)
  wire _00962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10573" *)
  wire _00963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10601" *)
  wire _00964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10621" *)
  wire _00965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10642" *)
  wire _00966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10650" *)
  wire _00967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10670" *)
  wire _00968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10670" *)
  wire _00969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10671" *)
  wire _00970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10672" *)
  wire _00971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10672" *)
  wire _00972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10673" *)
  wire _00973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10673" *)
  wire _00974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10681" *)
  wire _00975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10681" *)
  wire _00976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10690" *)
  wire _00977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10699" *)
  wire _00978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10707" *)
  wire _00979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10709" *)
  wire [31:0] _00980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10745" *)
  wire _00981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10745" *)
  wire _00982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10773" *)
  wire _00983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10781" *)
  wire _00984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10789" *)
  wire _00985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10790" *)
  wire _00986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10790" *)
  wire _00987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10799" *)
  wire _00988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10801" *)
  wire [31:0] _00989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10808" *)
  wire _00990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10808" *)
  wire _00991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10809" *)
  wire _00992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10809" *)
  wire _00993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10810" *)
  wire _00994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10810" *)
  wire _00995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10810" *)
  wire _00996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10818" *)
  wire _00997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10818" *)
  wire _00998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10819" *)
  wire _00999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10819" *)
  wire _01000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10828" *)
  wire _01001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10837" *)
  wire _01002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10845" *)
  wire _01003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10853" *)
  wire _01004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10874" *)
  wire _01005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10883" *)
  wire _01006_;
  wire [5:0] _01007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10893" *)
  wire _01008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10893" *)
  wire _01009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10901" *)
  wire _01010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10921" *)
  wire _01011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10922" *)
  wire _01012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10922" *)
  wire _01013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10931" *)
  wire _01014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10933" *)
  wire [31:0] _01015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10940" *)
  wire _01016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10940" *)
  wire _01017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10941" *)
  wire _01018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10941" *)
  wire _01019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10942" *)
  wire _01020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10942" *)
  wire _01021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10942" *)
  wire _01022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10950" *)
  wire _01023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10950" *)
  wire _01024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10951" *)
  wire _01025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10951" *)
  wire _01026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10960" *)
  wire _01027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10969" *)
  wire _01028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10977" *)
  wire _01029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10985" *)
  wire _01030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10994" *)
  wire _01031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11003" *)
  wire _01032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11005" *)
  wire [31:0] _01033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11013" *)
  wire _01034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11013" *)
  wire _01035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11021" *)
  wire _01036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11029" *)
  wire _01037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11030" *)
  wire _01038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11030" *)
  wire _01039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11039" *)
  wire _01040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11041" *)
  wire [31:0] _01041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11048" *)
  wire _01042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11048" *)
  wire _01043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11049" *)
  wire _01044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11049" *)
  wire _01045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11050" *)
  wire _01046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11050" *)
  wire _01047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11050" *)
  wire _01048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11058" *)
  wire _01049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11058" *)
  wire _01050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11059" *)
  wire _01051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11059" *)
  wire _01052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11068" *)
  wire _01053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11087" *)
  wire _01054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11095" *)
  wire _01055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11103" *)
  wire _01056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11111" *)
  wire _01057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11120" *)
  wire _01058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11129" *)
  wire _01059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11131" *)
  wire [31:0] _01060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11139" *)
  wire _01061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11139" *)
  wire _01062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11147" *)
  wire _01063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11155" *)
  wire _01064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11156" *)
  wire _01065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11156" *)
  wire _01066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11165" *)
  wire _01067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11167" *)
  wire [31:0] _01068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11174" *)
  wire _01069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11174" *)
  wire _01070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11175" *)
  wire _01071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11175" *)
  wire _01072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11176" *)
  wire _01073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11176" *)
  wire _01074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11176" *)
  wire _01075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11184" *)
  wire _01076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11184" *)
  wire _01077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11185" *)
  wire _01078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11185" *)
  wire _01079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11194" *)
  wire _01080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11218" *)
  wire _01081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11218" *)
  wire _01082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11227" *)
  wire _01083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11235" *)
  wire _01084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11243" *)
  wire _01085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11251" *)
  wire _01086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11271" *)
  wire _01087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11279" *)
  wire _01088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11287" *)
  wire _01089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11295" *)
  wire _01090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11303" *)
  wire _01091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11311" *)
  wire _01092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11329" *)
  wire _01093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11351" *)
  wire [7:0] _01094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11351" *)
  wire [7:0] _01095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11354" *)
  wire [7:0] _01096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11354" *)
  wire [7:0] _01097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11357" *)
  wire [7:0] _01098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11357" *)
  wire [7:0] _01099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11360" *)
  wire [7:0] _01100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11360" *)
  wire [7:0] _01101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11375" *)
  wire _01102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11375" *)
  wire _01103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11384" *)
  wire _01104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11392" *)
  wire _01105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11393" *)
  wire _01106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11402" *)
  wire _01107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11411" *)
  wire _01108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11420" *)
  wire _01109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11420" *)
  wire _01110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11429" *)
  wire _01111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11438" *)
  wire _01112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11457" *)
  wire _01113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11466" *)
  wire _01114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11475" *)
  wire _01115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11484" *)
  wire _01116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11504" *)
  wire _01117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11505" *)
  wire _01118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11515" *)
  wire _01119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11523" *)
  wire _01120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11533" *)
  wire _01121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11543" *)
  wire _01122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11551" *)
  wire _01123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11561" *)
  wire _01124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11571" *)
  wire _01125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11579" *)
  wire _01126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11589" *)
  wire _01127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11599" *)
  wire _01128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11607" *)
  wire _01129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11615" *)
  wire _01130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11623" *)
  wire _01131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11631" *)
  wire _01132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11649" *)
  wire _01133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11657" *)
  wire _01134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11665" *)
  wire _01135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11685" *)
  wire _01136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11747" *)
  wire [5:0] _01137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11750" *)
  wire [5:0] _01138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11753" *)
  wire [5:0] _01139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11756" *)
  wire [5:0] _01140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11759" *)
  wire _01141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11800" *)
  wire _01142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11841" *)
  wire _01143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11882" *)
  wire _01144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12040" *)
  wire _01145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12170" *)
  wire _01146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12235" *)
  wire _01147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12271" *)
  wire _01148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12271" *)
  wire _01149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12292" *)
  wire _01150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12298" *)
  wire _01151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12299" *)
  wire _01152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12313" *)
  wire _01153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12319" *)
  wire _01154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12320" *)
  wire _01155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12333" *)
  wire _01156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12339" *)
  wire _01157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12353" *)
  wire _01158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12360" *)
  wire _01159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12372" *)
  wire _01160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12419" *)
  wire _01161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12474" *)
  wire _01162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12517" *)
  wire _01163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12628" *)
  wire _01164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12637" *)
  wire _01165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12643" *)
  wire _01166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12652" *)
  wire _01167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12660" *)
  wire _01168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12660" *)
  wire _01169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12662" *)
  wire _01170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12667" *)
  wire _01171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12671" *)
  wire _01172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12671" *)
  wire _01173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12673" *)
  wire _01174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12678" *)
  wire _01175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12681" *)
  wire _01176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12681" *)
  wire _01177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12683" *)
  wire _01178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12688" *)
  wire _01179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12689" *)
  wire _01180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12720" *)
  wire _01181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12737" *)
  wire _01182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12754" *)
  wire _01183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12782" *)
  wire _01184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12792" *)
  wire _01185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12815" *)
  wire _01186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12815" *)
  wire _01187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12821" *)
  wire _01188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12821" *)
  wire _01189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12821" *)
  wire _01190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12822" *)
  wire _01191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12822" *)
  wire _01192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12852" *)
  wire _01193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12862" *)
  wire _01194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12862" *)
  wire _01195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12866" *)
  wire _01196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *)
  wire _01197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *)
  wire _01198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *)
  wire _01199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *)
  wire _01200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12870" *)
  wire _01201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12870" *)
  wire _01202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12871" *)
  wire _01203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12871" *)
  wire _01204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12871" *)
  wire _01205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12887" *)
  wire _01206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12899" *)
  wire _01207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12913" *)
  wire _01208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *)
  wire _01209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *)
  wire _01210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *)
  wire _01211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *)
  wire _01212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12917" *)
  wire _01213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12917" *)
  wire _01214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12918" *)
  wire _01215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12918" *)
  wire _01216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12918" *)
  wire _01217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12932" *)
  wire _01218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12939" *)
  wire _01219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12945" *)
  wire _01220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12955" *)
  wire _01221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12974" *)
  wire _01222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12974" *)
  wire _01223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12977" *)
  wire _01224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12977" *)
  wire _01225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12977" *)
  wire _01226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12978" *)
  wire _01227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12978" *)
  wire _01228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12982" *)
  wire _01229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12982" *)
  wire _01230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12993" *)
  wire _01231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12999" *)
  wire _01232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12999" *)
  wire _01233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13016" *)
  wire _01234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13016" *)
  wire _01235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13032" *)
  wire _01236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13032" *)
  wire _01237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13048" *)
  wire _01238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13048" *)
  wire _01239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13074" *)
  wire _01240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13079" *)
  wire _01241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13080" *)
  wire _01242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13115" *)
  wire _01243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13121" *)
  wire _01244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13122" *)
  wire _01245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13132" *)
  wire _01246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13134" *)
  wire _01247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13134" *)
  wire _01248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13136" *)
  wire _01249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13143" *)
  wire _01250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13143" *)
  wire _01251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13143" *)
  wire _01252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13144" *)
  wire _01253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13159" *)
  wire _01254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13160" *)
  wire _01255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13160" *)
  wire _01256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13164" *)
  wire _01257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13164" *)
  wire _01258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13176" *)
  wire _01259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13177" *)
  wire _01260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13177" *)
  wire _01261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13184" *)
  wire _01262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13186" *)
  wire _01263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13186" *)
  wire _01264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13188" *)
  wire _01265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13194" *)
  wire _01266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13195" *)
  wire _01267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13195" *)
  wire _01268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13198" *)
  wire _01269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13199" *)
  wire _01270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13201" *)
  wire _01271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13209" *)
  wire _01272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13209" *)
  wire _01273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13209" *)
  wire _01274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13211" *)
  wire _01275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13214" *)
  wire _01276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13216" *)
  wire _01277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13219" *)
  wire _01278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13221" *)
  wire _01279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13221" *)
  wire _01280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13234" *)
  wire _01281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13239" *)
  wire _01282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13247" *)
  wire _01283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13252" *)
  wire _01284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13260" *)
  wire _01285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13265" *)
  wire _01286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *)
  wire _01300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _01314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _01327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *)
  wire _01328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *)
  wire _01329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *)
  wire _01330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *)
  wire _01331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *)
  wire _01332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *)
  wire _01333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *)
  wire _01334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *)
  wire _01335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _01336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _01337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _01338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _01339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _01340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _01341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _01342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _01343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _01344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _01345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _01346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _01347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _01348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _01349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _01350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _01351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _01352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _01353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _01354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _01355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _01356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _01357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _01358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _01359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13318" *)
  wire [11:0] _01360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13318" *)
  wire [11:0] _01361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13318" *)
  wire [11:0] _01362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13318" *)
  wire [11:0] _01363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *)
  wire [11:0] _01364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *)
  wire [11:0] _01365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *)
  wire [11:0] _01366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *)
  wire [11:0] _01367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *)
  wire [11:0] _01368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *)
  wire [11:0] _01369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *)
  wire [11:0] _01370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *)
  wire [11:0] _01371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *)
  wire [11:0] _01372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *)
  wire [11:0] _01373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *)
  wire [11:0] _01374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *)
  wire [11:0] _01375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *)
  wire [11:0] _01376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *)
  wire [11:0] _01377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *)
  wire [11:0] _01378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *)
  wire [11:0] _01379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13336" *)
  wire [22:0] _01380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13336" *)
  wire [22:0] _01381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13336" *)
  wire [22:0] _01382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13336" *)
  wire [22:0] _01383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *)
  wire [22:0] _01384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *)
  wire [22:0] _01385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *)
  wire [22:0] _01386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *)
  wire [22:0] _01387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *)
  wire [22:0] _01388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *)
  wire [22:0] _01389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *)
  wire [22:0] _01390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *)
  wire [22:0] _01391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *)
  wire [22:0] _01392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *)
  wire [22:0] _01393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *)
  wire [22:0] _01394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *)
  wire [22:0] _01395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *)
  wire [22:0] _01396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *)
  wire [22:0] _01397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *)
  wire [22:0] _01398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *)
  wire [22:0] _01399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *)
  wire [22:0] _01400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *)
  wire [22:0] _01401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *)
  wire [22:0] _01402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *)
  wire [22:0] _01403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13352" *)
  wire [1:0] _01404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13352" *)
  wire [1:0] _01405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13352" *)
  wire [1:0] _01406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13352" *)
  wire [1:0] _01407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *)
  wire [1:0] _01408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *)
  wire [1:0] _01409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *)
  wire [1:0] _01410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *)
  wire [1:0] _01411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *)
  wire [1:0] _01412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *)
  wire [1:0] _01413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *)
  wire [1:0] _01414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *)
  wire [1:0] _01415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13366" *)
  wire [49:0] _01416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13366" *)
  wire [49:0] _01417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13366" *)
  wire [49:0] _01418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13366" *)
  wire [49:0] _01419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *)
  wire [49:0] _01420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *)
  wire [49:0] _01421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *)
  wire [49:0] _01422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *)
  wire [49:0] _01423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *)
  wire [49:0] _01424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *)
  wire [49:0] _01425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *)
  wire [49:0] _01426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *)
  wire [49:0] _01427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *)
  wire [49:0] _01428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *)
  wire [49:0] _01429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *)
  wire [49:0] _01430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *)
  wire [49:0] _01431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13380" *)
  wire [5:0] _01432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13380" *)
  wire [5:0] _01433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13380" *)
  wire [5:0] _01434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13380" *)
  wire [5:0] _01435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *)
  wire [5:0] _01436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *)
  wire [5:0] _01437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *)
  wire [5:0] _01438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *)
  wire [5:0] _01439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *)
  wire [5:0] _01440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *)
  wire [5:0] _01441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *)
  wire [5:0] _01442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *)
  wire [5:0] _01443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13396" *)
  wire [5:0] _01444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13396" *)
  wire [5:0] _01445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13396" *)
  wire [5:0] _01446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13396" *)
  wire [5:0] _01447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *)
  wire [5:0] _01448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *)
  wire [5:0] _01449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *)
  wire [5:0] _01450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *)
  wire [5:0] _01451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *)
  wire [5:0] _01452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *)
  wire [5:0] _01453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *)
  wire [5:0] _01454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *)
  wire [5:0] _01455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *)
  wire [5:0] _01456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *)
  wire [5:0] _01457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *)
  wire [5:0] _01458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *)
  wire [5:0] _01459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *)
  wire [5:0] _01460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *)
  wire [5:0] _01461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *)
  wire [5:0] _01462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *)
  wire [5:0] _01463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *)
  wire [5:0] _01464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *)
  wire [5:0] _01465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *)
  wire [5:0] _01466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *)
  wire [5:0] _01467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13412" *)
  wire [7:0] _01468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13412" *)
  wire [7:0] _01469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13412" *)
  wire [7:0] _01470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13412" *)
  wire [7:0] _01471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *)
  wire [7:0] _01472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *)
  wire [7:0] _01473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *)
  wire [7:0] _01474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *)
  wire [7:0] _01475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *)
  wire [7:0] _01476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *)
  wire [7:0] _01477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *)
  wire [7:0] _01478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *)
  wire [7:0] _01479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *)
  wire [7:0] _01480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *)
  wire [7:0] _01481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *)
  wire [7:0] _01482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *)
  wire [7:0] _01483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *)
  wire [7:0] _01484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *)
  wire [7:0] _01485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *)
  wire [7:0] _01486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *)
  wire [7:0] _01487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _01488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _01489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _01490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _01491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _01492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _01493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _01494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _01495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _01496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _01497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _01498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _01499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _01500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _01501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _01502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _01503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _01504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _01505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _01506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _01507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _01508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _01509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _01510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _01511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *)
  wire [7:0] _01512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *)
  wire [7:0] _01513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *)
  wire [7:0] _01514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *)
  wire [7:0] _01515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *)
  wire [7:0] _01516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *)
  wire [7:0] _01517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *)
  wire [7:0] _01518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *)
  wire [7:0] _01519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13444" *)
  wire [8:0] _01520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13444" *)
  wire [8:0] _01521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13444" *)
  wire [8:0] _01522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13444" *)
  wire [8:0] _01523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *)
  wire [8:0] _01524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *)
  wire [8:0] _01525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *)
  wire [8:0] _01526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *)
  wire [8:0] _01527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13446" *)
  wire [8:0] _01528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *)
  wire [8:0] _01529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *)
  wire [8:0] _01530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *)
  wire [8:0] _01531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *)
  wire [8:0] _01532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13448" *)
  wire [8:0] _01533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5453" *)
  wire _01534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5455" *)
  wire _01535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5457" *)
  wire _01536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5459" *)
  wire _01537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5483" *)
  wire _01538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5495" *)
  wire _01539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5527" *)
  wire _01540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5528" *)
  wire _01541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5551" *)
  wire _01542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5553" *)
  wire _01543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5559" *)
  wire _01544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5570" *)
  wire _01545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5572" *)
  wire _01546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5575" *)
  wire _01547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5577" *)
  wire _01548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5601" *)
  wire _01549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5603" *)
  wire _01550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5615" *)
  wire _01551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5617" *)
  wire _01552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5641" *)
  wire _01553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5643" *)
  wire _01554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5649" *)
  wire _01555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5651" *)
  wire _01556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5672" *)
  wire _01557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5674" *)
  wire _01558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5679" *)
  wire _01559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5681" *)
  wire _01560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5700" *)
  wire _01561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5776" *)
  wire _01562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5799" *)
  wire _01563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5803" *)
  wire _01564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5807" *)
  wire _01565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5809" *)
  wire _01566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5811" *)
  wire _01567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5813" *)
  wire _01568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5813" *)
  wire _01569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5814" *)
  wire _01570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5814" *)
  wire _01571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5814" *)
  wire _01572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5819" *)
  wire _01573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5821" *)
  wire _01574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5821" *)
  wire _01575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5823" *)
  wire _01576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5827" *)
  wire _01577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5829" *)
  wire _01578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5831" *)
  wire _01579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5834" *)
  wire _01580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5836" *)
  wire _01581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5841" *)
  wire _01582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5841" *)
  wire _01583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5843" *)
  wire _01584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5844" *)
  wire _01585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5846" *)
  wire _01586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5852" *)
  wire _01587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5853" *)
  wire _01588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5854" *)
  wire _01589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5855" *)
  wire _01590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5857" *)
  wire _01591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5857" *)
  wire _01592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5860" *)
  wire _01593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5861" *)
  wire _01594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5865" *)
  wire _01595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5871" *)
  wire _01596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5887" *)
  wire _01597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5887" *)
  wire _01598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5894" *)
  wire _01599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5895" *)
  wire _01600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5896" *)
  wire _01601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5897" *)
  wire _01602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5902" *)
  wire _01603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5903" *)
  wire _01604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5982" *)
  wire _01605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5989" *)
  wire _01606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5991" *)
  wire _01607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5996" *)
  wire _01608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6014" *)
  wire _01609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6040" *)
  wire _01610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6048" *)
  wire _01611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6060" *)
  wire _01612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6092" *)
  wire _01613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6133" *)
  wire _01614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6598" *)
  wire _01615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6626" *)
  wire _01616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6649" *)
  wire _01617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6679" *)
  wire _01618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6702" *)
  wire _01619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6730" *)
  wire _01620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6753" *)
  wire _01621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6781" *)
  wire _01622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6871" *)
  wire [34:0] _01623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6871" *)
  wire [34:0] _01624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6872" *)
  wire [34:0] _01625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6889" *)
  wire [7:0] _01626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6894" *)
  wire [34:0] _01627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6894" *)
  wire [34:0] _01628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6895" *)
  wire [34:0] _01629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6929" *)
  wire [34:0] _01630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6929" *)
  wire [34:0] _01631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6930" *)
  wire [34:0] _01632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6947" *)
  wire [7:0] _01633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6952" *)
  wire [34:0] _01634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6952" *)
  wire [34:0] _01635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6953" *)
  wire [34:0] _01636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6987" *)
  wire [34:0] _01637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6987" *)
  wire [34:0] _01638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6988" *)
  wire [34:0] _01639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7005" *)
  wire [7:0] _01640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7010" *)
  wire [34:0] _01641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7010" *)
  wire [34:0] _01642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7011" *)
  wire [34:0] _01643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7045" *)
  wire [34:0] _01644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7045" *)
  wire [34:0] _01645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7046" *)
  wire [34:0] _01646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7063" *)
  wire [7:0] _01647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7068" *)
  wire [34:0] _01648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7068" *)
  wire [34:0] _01649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7069" *)
  wire [34:0] _01650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7075" *)
  wire _01651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7077" *)
  wire _01652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7079" *)
  wire _01653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7081" *)
  wire _01654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7083" *)
  wire _01655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7084" *)
  wire _01656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7085" *)
  wire _01657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7085" *)
  wire _01658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7085" *)
  wire _01659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7091" *)
  wire _01660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7093" *)
  wire _01661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7095" *)
  wire _01662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7097" *)
  wire _01663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7098" *)
  wire _01664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7099" *)
  wire _01665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7099" *)
  wire _01666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7099" *)
  wire _01667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7109" *)
  wire _01668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7111" *)
  wire _01669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7112" *)
  wire _01670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7113" *)
  wire _01671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7113" *)
  wire _01672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7113" *)
  wire _01673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7123" *)
  wire _01674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7125" *)
  wire _01675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7126" *)
  wire _01676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7127" *)
  wire _01677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7127" *)
  wire _01678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7127" *)
  wire _01679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7468" *)
  wire _01680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7478" *)
  wire _01681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7482" *)
  wire _01682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7487" *)
  wire _01683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7490" *)
  wire _01684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7498" *)
  wire _01685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7509" *)
  wire _01686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7509" *)
  wire _01687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7515" *)
  wire _01688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7517" *)
  wire _01689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7519" *)
  wire _01690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7528" *)
  wire _01691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7529" *)
  wire _01692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7533" *)
  wire _01693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7534" *)
  wire _01694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7535" *)
  wire _01695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7538" *)
  wire _01696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7539" *)
  wire _01697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7541" *)
  wire _01698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7545" *)
  wire _01699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7546" *)
  wire _01700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7552" *)
  wire _01701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7561" *)
  wire _01702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7561" *)
  wire _01703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7565" *)
  wire _01704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7571" *)
  wire _01705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7576" *)
  wire _01706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7604" *)
  wire _01707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7611" *)
  wire _01708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7612" *)
  wire _01709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7615" *)
  wire _01710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7625" *)
  wire _01711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7625" *)
  wire _01712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7625" *)
  wire _01713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7626" *)
  wire _01714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7626" *)
  wire _01715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7628" *)
  wire _01716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7628" *)
  wire _01717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7631" *)
  wire _01718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7635" *)
  wire _01719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7635" *)
  wire _01720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7637" *)
  wire _01721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7637" *)
  wire _01722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7637" *)
  wire _01723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7638" *)
  wire _01724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7638" *)
  wire _01725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7640" *)
  wire _01726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7640" *)
  wire _01727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *)
  wire _01728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *)
  wire _01729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7644" *)
  wire _01730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7644" *)
  wire _01731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7646" *)
  wire _01732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7646" *)
  wire _01733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7646" *)
  wire _01734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7647" *)
  wire _01735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7647" *)
  wire _01736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7649" *)
  wire _01737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7649" *)
  wire _01738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7652" *)
  wire _01739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7654" *)
  wire _01740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7654" *)
  wire _01741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7656" *)
  wire _01742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7656" *)
  wire _01743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7656" *)
  wire _01744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7657" *)
  wire _01745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7657" *)
  wire _01746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7663" *)
  wire _01747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7663" *)
  wire _01748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7667" *)
  wire _01749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7667" *)
  wire _01750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7680" *)
  wire _01751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7722" *)
  wire _01752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7725" *)
  wire _01753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7727" *)
  wire _01754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7729" *)
  wire _01755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7731" *)
  wire _01756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7733" *)
  wire _01757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7734" *)
  wire _01758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7737" *)
  wire _01759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7744" *)
  wire _01760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7745" *)
  wire _01761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7748" *)
  wire _01762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7749" *)
  wire _01763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7750" *)
  wire _01764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7751" *)
  wire _01765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7752" *)
  wire _01766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7754" *)
  wire _01767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7759" *)
  wire _01768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7764" *)
  wire _01769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7769" *)
  wire _01770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7813" *)
  wire _01771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7816" *)
  wire _01772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7886" *)
  wire _01773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7894" *)
  wire _01774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7960" *)
  wire _01775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7961" *)
  wire _01776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7962" *)
  wire _01777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7963" *)
  wire _01778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8086" *)
  wire _01779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8094" *)
  wire _01780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8139" *)
  wire _01781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8224" *)
  wire _01782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8224" *)
  wire _01783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8268" *)
  wire _01784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8269" *)
  wire _01785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8269" *)
  wire _01786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8278" *)
  wire _01787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8278" *)
  wire _01788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8278" *)
  wire _01789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8287" *)
  wire _01790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8287" *)
  wire _01791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8310" *)
  wire _01792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8311" *)
  wire _01793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8311" *)
  wire _01794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8333" *)
  wire _01795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8333" *)
  wire _01796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8333" *)
  wire _01797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8342" *)
  wire _01798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8342" *)
  wire _01799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8363" *)
  wire _01800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8364" *)
  wire _01801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8364" *)
  wire _01802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8373" *)
  wire _01803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8374" *)
  wire _01804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8374" *)
  wire _01805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8383" *)
  wire _01806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8383" *)
  wire _01807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8412" *)
  wire _01808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8413" *)
  wire _01809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8413" *)
  wire _01810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8422" *)
  wire _01811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8423" *)
  wire _01812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8423" *)
  wire _01813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8432" *)
  wire _01814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8432" *)
  wire _01815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8443" *)
  wire _01816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8444" *)
  wire _01817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8444" *)
  wire _01818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8453" *)
  wire _01819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8453" *)
  wire _01820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8503" *)
  wire _01821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8504" *)
  wire _01822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8515" *)
  wire _01823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8525" *)
  wire _01824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8525" *)
  wire _01825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8526" *)
  wire _01826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8526" *)
  wire _01827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8547" *)
  wire _01828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8548" *)
  wire _01829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8548" *)
  wire _01830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8558" *)
  wire _01831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8558" *)
  wire _01832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8568" *)
  wire _01833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8568" *)
  wire _01834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8645" *)
  wire _01835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8655" *)
  wire _01836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8665" *)
  wire _01837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8676" *)
  wire _01838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8676" *)
  wire _01839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8687" *)
  wire _01840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8696" *)
  wire _01841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8723" *)
  wire _01842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8724" *)
  wire _01843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8735" *)
  wire _01844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8745" *)
  wire _01845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8745" *)
  wire _01846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8746" *)
  wire _01847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8746" *)
  wire _01848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8768" *)
  wire _01849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8768" *)
  wire _01850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8768" *)
  wire _01851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8778" *)
  wire _01852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8778" *)
  wire _01853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8788" *)
  wire _01854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8814" *)
  wire _01855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8824" *)
  wire _01856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8835" *)
  wire _01857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8836" *)
  wire _01858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8862" *)
  wire _01859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8872" *)
  wire _01860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8883" *)
  wire _01861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8893" *)
  wire _01862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8893" *)
  wire _01863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8894" *)
  wire _01864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8894" *)
  wire _01865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8916" *)
  wire _01866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8917" *)
  wire _01867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8917" *)
  wire _01868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8927" *)
  wire _01869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8927" *)
  wire _01870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8937" *)
  wire _01871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8948" *)
  wire _01872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8958" *)
  wire _01873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8969" *)
  wire _01874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8970" *)
  wire _01875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8982" *)
  wire _01876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8992" *)
  wire _01877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9003" *)
  wire _01878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9013" *)
  wire _01879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9013" *)
  wire _01880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9014" *)
  wire _01881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9014" *)
  wire _01882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9036" *)
  wire _01883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9037" *)
  wire _01884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9037" *)
  wire _01885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9047" *)
  wire _01886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9047" *)
  wire _01887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9057" *)
  wire _01888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9068" *)
  wire _01889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9078" *)
  wire _01890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9089" *)
  wire _01891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9090" *)
  wire _01892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9102" *)
  wire _01893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9111" *)
  wire _01894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9111" *)
  wire _01895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9129" *)
  wire _01896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9139" *)
  wire _01897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9185" *)
  wire [5:0] _01898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9185" *)
  wire [5:0] _01899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9186" *)
  wire [5:0] _01900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9191" *)
  wire [5:0] _01901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9191" *)
  wire [5:0] _01902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9192" *)
  wire [5:0] _01903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9197" *)
  wire [5:0] _01904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9197" *)
  wire [5:0] _01905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9198" *)
  wire [5:0] _01906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9203" *)
  wire [5:0] _01907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9203" *)
  wire [5:0] _01908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9204" *)
  wire [5:0] _01909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9223" *)
  wire _01910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9224" *)
  wire _01911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9244" *)
  wire _01912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9255" *)
  wire _01913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9265" *)
  wire _01914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9284" *)
  wire _01915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9304" *)
  wire _01916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9315" *)
  wire _01917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9325" *)
  wire _01918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9344" *)
  wire _01919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9364" *)
  wire _01920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9375" *)
  wire _01921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9385" *)
  wire _01922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9404" *)
  wire _01923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9424" *)
  wire _01924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9433" *)
  wire _01925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9433" *)
  wire _01926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9490" *)
  wire [22:0] _01927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9490" *)
  wire [22:0] _01928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9491" *)
  wire [22:0] _01929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9494" *)
  wire [34:0] _01930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9494" *)
  wire [34:0] _01931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9495" *)
  wire [34:0] _01932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9498" *)
  wire [34:0] _01933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9498" *)
  wire [34:0] _01934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9501" *)
  wire [34:0] _01935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9501" *)
  wire [34:0] _01936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9505" *)
  wire [22:0] _01937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9505" *)
  wire [22:0] _01938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9506" *)
  wire [22:0] _01939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9509" *)
  wire [34:0] _01940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9509" *)
  wire [34:0] _01941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9510" *)
  wire [34:0] _01942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9513" *)
  wire [34:0] _01943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9513" *)
  wire [34:0] _01944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9516" *)
  wire [34:0] _01945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9516" *)
  wire [34:0] _01946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9519" *)
  wire [22:0] _01947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9519" *)
  wire [22:0] _01948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9520" *)
  wire [22:0] _01949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9523" *)
  wire [34:0] _01950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9523" *)
  wire [34:0] _01951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9524" *)
  wire [34:0] _01952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9527" *)
  wire [34:0] _01953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9527" *)
  wire [34:0] _01954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9530" *)
  wire [34:0] _01955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9530" *)
  wire [34:0] _01956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9533" *)
  wire [22:0] _01957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9533" *)
  wire [22:0] _01958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9534" *)
  wire [22:0] _01959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9537" *)
  wire [34:0] _01960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9537" *)
  wire [34:0] _01961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9538" *)
  wire [34:0] _01962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9541" *)
  wire [34:0] _01963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9541" *)
  wire [34:0] _01964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9544" *)
  wire [34:0] _01965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9544" *)
  wire [34:0] _01966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9546" *)
  wire _01967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9547" *)
  wire _01968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9548" *)
  wire _01969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9550" *)
  wire _01970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9553" *)
  wire [5:0] _01971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9553" *)
  wire [5:0] _01972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9554" *)
  wire [5:0] _01973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9562" *)
  wire [5:0] _01974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9562" *)
  wire [5:0] _01975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9563" *)
  wire [5:0] _01976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9568" *)
  wire [5:0] _01977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9568" *)
  wire [5:0] _01978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9569" *)
  wire [5:0] _01979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9574" *)
  wire [5:0] _01980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9574" *)
  wire [5:0] _01981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9575" *)
  wire [5:0] _01982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9589" *)
  wire _01983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9590" *)
  wire _01984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9599" *)
  wire _01985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9608" *)
  wire _01986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9617" *)
  wire _01987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9625" *)
  wire _01988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9633" *)
  wire _01989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9653" *)
  wire _01990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9661" *)
  wire _01991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9670" *)
  wire _01992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9679" *)
  wire _01993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9687" *)
  wire _01994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9719" *)
  wire _01995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9720" *)
  wire _01996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9729" *)
  wire _01997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9738" *)
  wire _01998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9747" *)
  wire _01999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9755" *)
  wire _02000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9763" *)
  wire _02001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9771" *)
  wire _02002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9779" *)
  wire _02003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9788" *)
  wire _02004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9797" *)
  wire _02005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9805" *)
  wire _02006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9813" *)
  wire _02007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9814" *)
  wire _02008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9823" *)
  wire _02009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9832" *)
  wire _02010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9841" *)
  wire _02011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9849" *)
  wire _02012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9867" *)
  wire _02013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9876" *)
  wire _02014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9885" *)
  wire _02015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9893" *)
  wire _02016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9911" *)
  wire _02017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9912" *)
  wire _02018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9921" *)
  wire _02019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9930" *)
  wire _02020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9939" *)
  wire _02021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9947" *)
  wire _02022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9955" *)
  wire _02023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9964" *)
  wire _02024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9973" *)
  wire _02025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9981" *)
  wire _02026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10885" *)
  wire [31:0] _02027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7055" *)
  wire [246:0] _02028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4444" *)
  wire [7:0] _02029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4286" *)
  (* unused_bits = "9" *)
  wire [9:0] _02030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13078" *)
  wire _02031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13120" *)
  wire _02032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5962" *)
  wire _02033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6010" *)
  wire _02034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6057" *)
  wire _02035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6097" *)
  wire _02036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6138" *)
  wire _02037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6153" *)
  wire _02038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6154" *)
  wire _02039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6155" *)
  wire _02040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6156" *)
  wire _02041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6216" *)
  wire _02042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6232" *)
  wire _02043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6256" *)
  wire _02044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6272" *)
  wire _02045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6296" *)
  wire _02046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6312" *)
  wire _02047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6336" *)
  wire _02048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6352" *)
  wire _02049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6414" *)
  wire _02050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6475" *)
  wire _02051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6481" *)
  wire _02052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6662" *)
  wire _02053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7541" *)
  wire _02054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10222" *)
  wire _02055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12380" *)
  wire _02056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12405" *)
  wire _02057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5961" *)
  wire _02058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5964" *)
  wire _02059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6009" *)
  wire _02060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6056" *)
  wire _02061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6096" *)
  wire _02062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6137" *)
  wire _02063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6191" *)
  wire _02064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6192" *)
  wire _02065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6368" *)
  wire _02066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6381" *)
  wire _02067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6396" *)
  wire _02068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6411" *)
  wire _02069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6474" *)
  wire _02070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6477" *)
  wire _02071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6480" *)
  wire _02072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6483" *)
  wire _02073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6485" *)
  wire _02074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6486" *)
  wire _02075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6550" *)
  wire _02076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6552" *)
  wire _02077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7325" *)
  wire _02078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7326" *)
  wire _02079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7331" *)
  wire _02080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7336" *)
  wire _02081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7379" *)
  wire _02082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7385" *)
  wire _02083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7391" *)
  wire _02084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7397" *)
  wire _02085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7403" *)
  wire _02086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7409" *)
  wire _02087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7415" *)
  wire _02088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7421" *)
  wire _02089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7456" *)
  wire _02090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7458" *)
  wire _02091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7460" *)
  wire _02092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7462" *)
  wire _02093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8197" *)
  wire _02094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8211" *)
  wire _02095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10072" *)
  wire _02096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10074" *)
  wire _02097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10076" *)
  wire _02098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10078" *)
  wire _02099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10108" *)
  wire _02100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10204" *)
  wire _02101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10204" *)
  wire _02102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10230" *)
  wire _02103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10310" *)
  wire _02104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10319" *)
  wire _02105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10321" *)
  wire _02106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10330" *)
  wire _02107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10341" *)
  wire _02108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10363" *)
  wire _02109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10385" *)
  wire _02110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10526" *)
  wire _02111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10670" *)
  wire _02112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10671" *)
  wire _02113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10673" *)
  wire _02114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10744" *)
  wire _02115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10790" *)
  wire _02116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10799" *)
  wire _02117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10808" *)
  wire _02118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10809" *)
  wire _02119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10818" *)
  wire _02120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10892" *)
  wire _02121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10922" *)
  wire _02122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10931" *)
  wire _02123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10940" *)
  wire _02124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10941" *)
  wire _02125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10950" *)
  wire _02126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11012" *)
  wire _02127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11030" *)
  wire _02128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11039" *)
  wire _02129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11048" *)
  wire _02130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11049" *)
  wire _02131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11138" *)
  wire _02132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11156" *)
  wire _02133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11165" *)
  wire _02134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11174" *)
  wire _02135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11175" *)
  wire _02136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11206" *)
  wire _02137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11208" *)
  wire _02138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11210" *)
  wire _02139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11219" *)
  wire _02140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11350" *)
  wire _02141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11353" *)
  wire _02142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11356" *)
  wire _02143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11359" *)
  wire _02144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11377" *)
  wire _02145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11404" *)
  wire _02146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11523" *)
  wire _02147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11551" *)
  wire _02148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11579" *)
  wire _02149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11607" *)
  wire _02150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11615" *)
  wire _02151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11759" *)
  wire _02152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11800" *)
  wire _02153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11841" *)
  wire _02154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11882" *)
  wire _02155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11949" *)
  wire [48:0] _02156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11955" *)
  wire [48:0] _02157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11964" *)
  wire [48:0] _02158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11967" *)
  wire [48:0] _02159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11973" *)
  wire [48:0] _02160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11982" *)
  wire [48:0] _02161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11985" *)
  wire [48:0] _02162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11991" *)
  wire [48:0] _02163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12000" *)
  wire [48:0] _02164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12003" *)
  wire [48:0] _02165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12009" *)
  wire [48:0] _02166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12018" *)
  wire [48:0] _02167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12028" *)
  wire _02168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12031" *)
  wire _02169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12038" *)
  wire _02170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12040" *)
  wire _02171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12066" *)
  wire [5:0] _02172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12091" *)
  wire _02173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12098" *)
  wire _02174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12101" *)
  wire _02175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12107" *)
  wire _02176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12134" *)
  wire [5:0] _02177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12144" *)
  wire _02178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12157" *)
  wire _02179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12160" *)
  wire _02180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12170" *)
  wire _02181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12196" *)
  wire [5:0] _02182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12222" *)
  wire _02183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12225" *)
  wire _02184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12235" *)
  wire _02185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12262" *)
  wire [5:0] _02186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12273" *)
  wire _02187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12274" *)
  wire _02188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12280" *)
  wire _02189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12281" *)
  wire _02190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12283" *)
  wire _02191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12301" *)
  wire _02192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12302" *)
  wire _02193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12304" *)
  wire _02194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12322" *)
  wire _02195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12323" *)
  wire _02196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12341" *)
  wire _02197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12342" *)
  wire _02198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12344" *)
  wire _02199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12374" *)
  wire _02200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12375" *)
  wire _02201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12378" *)
  wire _02202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12380" *)
  wire _02203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12400" *)
  wire _02204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12403" *)
  wire _02205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12421" *)
  wire _02206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12425" *)
  wire _02207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12437" *)
  wire _02208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12457" *)
  wire _02209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12460" *)
  wire _02210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12476" *)
  wire _02211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12480" *)
  wire _02212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12498" *)
  wire _02213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12501" *)
  wire _02214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12519" *)
  wire _02215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12523" *)
  wire _02216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12541" *)
  wire _02217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12544" *)
  wire _02218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12557" *)
  wire _02219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12560" *)
  wire _02220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12563" *)
  wire _02221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12566" *)
  wire _02222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12569" *)
  wire _02223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12572" *)
  wire _02224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12575" *)
  wire _02225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12578" *)
  wire _02226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12612" *)
  wire _02227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12621" *)
  wire _02228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12622" *)
  wire _02229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12628" *)
  wire _02230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12643" *)
  wire _02231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12651" *)
  wire _02232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12692" *)
  wire _02233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12699" *)
  wire _02234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12701" *)
  wire _02235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12704" *)
  wire _02236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12705" *)
  wire _02237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12706" *)
  wire _02238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12713" *)
  wire _02239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12723" *)
  wire _02240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12724" *)
  wire _02241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12730" *)
  wire _02242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12740" *)
  wire _02243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12741" *)
  wire _02244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12746" *)
  wire _02245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12753" *)
  wire _02246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12754" *)
  wire _02247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12757" *)
  wire _02248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12758" *)
  wire _02249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12764" *)
  wire _02250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12768" *)
  wire _02251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12782" *)
  wire _02252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12810" *)
  wire _02253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12811" *)
  wire _02254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12815" *)
  wire _02255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12824" *)
  wire _02256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12833" *)
  wire _02257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12835" *)
  wire _02258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12837" *)
  wire _02259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12862" *)
  wire _02260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *)
  wire _02261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12873" *)
  wire _02262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12880" *)
  wire _02263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12882" *)
  wire _02264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12910" *)
  wire _02265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *)
  wire _02266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12920" *)
  wire _02267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12927" *)
  wire _02268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12929" *)
  wire _02269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12939" *)
  wire _02270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12945" *)
  wire _02271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12971" *)
  wire _02272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12974" *)
  wire _02273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12988" *)
  wire _02274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12990" *)
  wire _02275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12999" *)
  wire _02276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13016" *)
  wire _02277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13032" *)
  wire _02278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13048" *)
  wire _02279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13065" *)
  wire _02280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13066" *)
  wire _02281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13069" *)
  wire _02282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13074" *)
  wire _02283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13111" *)
  wire _02284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13115" *)
  wire _02285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13133" *)
  wire _02286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13134" *)
  wire _02287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13146" *)
  wire _02288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13147" *)
  wire _02289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13153" *)
  wire _02290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13164" *)
  wire _02291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13170" *)
  wire _02292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13179" *)
  wire _02293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13180" *)
  wire _02294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13185" *)
  wire _02295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13186" *)
  wire _02296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13199" *)
  wire _02297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13209" *)
  wire _02298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13211" *)
  wire _02299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13213" *)
  wire _02300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13214" *)
  wire _02301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13218" *)
  wire _02302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13219" *)
  wire _02303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13221" *)
  wire _02304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13236" *)
  wire _02305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13249" *)
  wire _02306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13262" *)
  wire _02307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13273" *)
  wire _02308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13276" *)
  wire _02309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4447" *)
  wire [6:0] _02310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4458" *)
  wire [6:0] _02311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4493" *)
  wire [6:0] _02312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4504" *)
  wire [6:0] _02313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4539" *)
  wire [6:0] _02314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4550" *)
  wire [6:0] _02315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4585" *)
  wire [6:0] _02316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4596" *)
  wire [6:0] _02317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5452" *)
  wire _02318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5461" *)
  wire _02319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5471" *)
  wire _02320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5483" *)
  wire _02321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5488" *)
  wire _02322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5496" *)
  wire _02323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5501" *)
  wire _02324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5503" *)
  wire _02325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5505" *)
  wire _02326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5510" *)
  wire _02327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5512" *)
  wire _02328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5519" *)
  wire _02329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5540" *)
  wire _02330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5542" *)
  wire [5:0] _02331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5550" *)
  wire _02332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5556" *)
  wire _02333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5562" *)
  wire _02334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5564" *)
  wire _02335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5569" *)
  wire _02336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5590" *)
  wire _02337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5592" *)
  wire [5:0] _02338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5600" *)
  wire _02339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5611" *)
  wire _02340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5614" *)
  wire _02341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5619" *)
  wire _02342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5620" *)
  wire _02343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5630" *)
  wire _02344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5632" *)
  wire [5:0] _02345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5640" *)
  wire _02346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5644" *)
  wire _02347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5648" *)
  wire _02348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5661" *)
  wire _02349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5663" *)
  wire [5:0] _02350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5671" *)
  wire _02351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5675" *)
  wire _02352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5678" *)
  wire _02353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5687" *)
  wire _02354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5688" *)
  wire _02355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5705" *)
  wire _02356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5717" *)
  wire _02357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5729" *)
  wire _02358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5740" *)
  wire _02359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5747" *)
  wire _02360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5754" *)
  wire _02361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5756" *)
  wire _02362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5768" *)
  wire _02363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5772" *)
  wire _02364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5780" *)
  wire _02365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5801" *)
  wire _02366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5810" *)
  wire _02367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5813" *)
  wire _02368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5818" *)
  wire _02369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5822" *)
  wire _02370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5826" *)
  wire _02371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5828" *)
  wire _02372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5830" *)
  wire _02373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5833" *)
  wire _02374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5835" *)
  wire _02375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5852" *)
  wire _02376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5853" *)
  wire _02377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5856" *)
  wire _02378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5862" *)
  wire _02379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5867" *)
  wire _02380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5869" *)
  wire _02381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5878" *)
  wire _02382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5884" *)
  wire _02383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5894" *)
  wire _02384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5895" *)
  wire _02385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5898" *)
  wire _02386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5900" *)
  wire _02387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5910" *)
  wire _02388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5912" *)
  wire _02389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5921" *)
  wire _02390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5925" *)
  wire _02391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5935" *)
  wire _02392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5956" *)
  wire _02393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5963" *)
  wire _02394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5982" *)
  wire _02395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6000" *)
  wire _02396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6014" *)
  wire _02397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6020" *)
  wire _02398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6040" *)
  wire _02399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6055" *)
  wire _02400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6060" *)
  wire _02401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6066" *)
  wire _02402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6084" *)
  wire _02403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6095" *)
  wire _02404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6108" *)
  wire _02405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6136" *)
  wire _02406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6416" *)
  wire _02407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6422" *)
  wire _02408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6428" *)
  wire _02409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6434" *)
  wire _02410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6476" *)
  wire _02411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6477" *)
  wire _02412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6482" *)
  wire _02413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6483" *)
  wire _02414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6485" *)
  wire _02415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6486" *)
  wire _02416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6587" *)
  wire _02417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6595" *)
  wire _02418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6597" *)
  wire _02419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6615" *)
  wire _02420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6623" *)
  wire _02421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6625" *)
  wire _02422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6638" *)
  wire _02423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6646" *)
  wire _02424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6648" *)
  wire _02425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6668" *)
  wire _02426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6676" *)
  wire _02427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6678" *)
  wire _02428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6691" *)
  wire _02429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6699" *)
  wire _02430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6701" *)
  wire _02431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6719" *)
  wire _02432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6727" *)
  wire _02433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6729" *)
  wire _02434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6742" *)
  wire _02435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6750" *)
  wire _02436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6752" *)
  wire _02437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6770" *)
  wire _02438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6778" *)
  wire _02439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6780" *)
  wire _02440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6874" *)
  wire [246:0] _02441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6881" *)
  wire [246:0] _02442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6932" *)
  wire [246:0] _02443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6939" *)
  wire [246:0] _02444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6990" *)
  wire [246:0] _02445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6997" *)
  wire [246:0] _02446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7048" *)
  wire [246:0] _02447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7075" *)
  wire _02448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7081" *)
  wire _02449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7084" *)
  wire _02450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7085" *)
  wire _02451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7089" *)
  wire _02452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7090" *)
  wire _02453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7095" *)
  wire _02454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7098" *)
  wire _02455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7099" *)
  wire _02456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7103" *)
  wire _02457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7109" *)
  wire _02458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7112" *)
  wire _02459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7113" *)
  wire _02460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7117" *)
  wire _02461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7123" *)
  wire _02462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7126" *)
  wire _02463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7127" *)
  wire _02464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7375" *)
  wire [1:0] _02465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7376" *)
  wire [5:0] _02466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7381" *)
  wire [7:0] _02467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7387" *)
  wire [1:0] _02468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7388" *)
  wire [5:0] _02469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7393" *)
  wire [7:0] _02470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7399" *)
  wire [1:0] _02471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7400" *)
  wire [5:0] _02472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7405" *)
  wire [7:0] _02473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7411" *)
  wire [1:0] _02474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7412" *)
  wire [5:0] _02475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7417" *)
  wire [7:0] _02476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7468" *)
  wire _02477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7478" *)
  wire _02478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7490" *)
  wire _02479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7498" *)
  wire _02480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7511" *)
  wire _02481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7584" *)
  wire _02482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7597" *)
  wire _02483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7604" *)
  wire _02484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7633" *)
  wire _02485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *)
  wire _02486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *)
  wire _02487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7652" *)
  wire _02488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7661" *)
  wire _02489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7674" *)
  wire _02490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7689" *)
  wire _02491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7690" *)
  wire _02492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7696" *)
  wire _02493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7697" *)
  wire _02494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7704" *)
  wire _02495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7705" *)
  wire _02496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7712" *)
  wire _02497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7713" *)
  wire _02498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7722" *)
  wire _02499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7723" *)
  wire _02500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7724" *)
  wire _02501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7725" *)
  wire _02502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7726" *)
  wire _02503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7727" *)
  wire _02504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7728" *)
  wire _02505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7729" *)
  wire _02506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7730" *)
  wire _02507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7731" *)
  wire _02508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7732" *)
  wire _02509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7733" *)
  wire _02510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7734" *)
  wire _02511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7735" *)
  wire _02512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7736" *)
  wire _02513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7737" *)
  wire _02514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7742" *)
  wire _02515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7754" *)
  wire _02516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7759" *)
  wire _02517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7764" *)
  wire _02518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7769" *)
  wire _02519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7789" *)
  wire [6:0] _02520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7792" *)
  wire [6:0] _02521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7795" *)
  wire [6:0] _02522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7798" *)
  wire [6:0] _02523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7801" *)
  wire [6:0] _02524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7804" *)
  wire [6:0] _02525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7807" *)
  wire [6:0] _02526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7810" *)
  wire [6:0] _02527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7814" *)
  wire _02528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7817" *)
  wire _02529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7823" *)
  wire _02530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7836" *)
  wire _02531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7838" *)
  wire _02532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7843" *)
  wire _02533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7851" *)
  wire _02534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7856" *)
  wire _02535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7860" *)
  wire _02536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7886" *)
  wire _02537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7988" *)
  wire _02538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7989" *)
  wire _02539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7990" *)
  wire _02540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7991" *)
  wire _02541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7992" *)
  wire _02542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7993" *)
  wire _02543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7994" *)
  wire _02544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7995" *)
  wire _02545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8087" *)
  wire _02546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8095" *)
  wire _02547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8197" *)
  wire _02548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8211" *)
  wire _02549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8217" *)
  wire _02550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8225" *)
  wire _02551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8310" *)
  wire _02552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8363" *)
  wire _02553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8412" *)
  wire _02554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8443" *)
  wire _02555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8454" *)
  wire _02556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8503" *)
  wire _02557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8515" *)
  wire _02558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8526" *)
  wire _02559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8558" *)
  wire _02560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8676" *)
  wire _02561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8687" *)
  wire _02562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8724" *)
  wire _02563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8735" *)
  wire _02564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8746" *)
  wire _02565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8778" *)
  wire _02566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8835" *)
  wire _02567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8872" *)
  wire _02568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8883" *)
  wire _02569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8894" *)
  wire _02570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8915" *)
  wire _02571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8927" *)
  wire _02572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8969" *)
  wire _02573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8992" *)
  wire _02574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9003" *)
  wire _02575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9014" *)
  wire _02576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9035" *)
  wire _02577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9047" *)
  wire _02578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9089" *)
  wire _02579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9112" *)
  wire _02580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9129" *)
  wire _02581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9185" *)
  wire _02582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9191" *)
  wire _02583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9197" *)
  wire _02584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9215" *)
  wire _02585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9235" *)
  wire _02586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9255" *)
  wire _02587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9315" *)
  wire _02588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9375" *)
  wire _02589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9434" *)
  wire _02590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9491" *)
  wire _02591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9494" *)
  wire _02592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9500" *)
  wire _02593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9506" *)
  wire _02594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9509" *)
  wire _02595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9515" *)
  wire _02596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9520" *)
  wire _02597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9523" *)
  wire _02598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9529" *)
  wire _02599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9534" *)
  wire _02600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9537" *)
  wire _02601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9543" *)
  wire _02602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9617" *)
  wire _02603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9633" *)
  wire _02604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9687" *)
  wire _02605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9763" *)
  wire _02606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9771" *)
  wire _02607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9797" *)
  wire _02608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9805" *)
  wire _02609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9841" *)
  wire _02610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9876" *)
  wire _02611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9885" *)
  wire _02612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9893" *)
  wire _02613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9939" *)
  wire _02614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9964" *)
  wire _02615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9973" *)
  wire _02616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9981" *)
  wire _02617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10307" *)
  wire _02618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10307" *)
  wire _02619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10318" *)
  wire _02620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10319" *)
  wire _02621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10319" *)
  wire _02622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10329" *)
  wire _02623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10329" *)
  wire _02624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10340" *)
  wire _02625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10341" *)
  wire _02626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10341" *)
  wire _02627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10351" *)
  wire _02628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10351" *)
  wire _02629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10362" *)
  wire _02630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10363" *)
  wire _02631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10363" *)
  wire _02632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10373" *)
  wire _02633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10373" *)
  wire _02634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10384" *)
  wire _02635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10385" *)
  wire _02636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10385" *)
  wire _02637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10673" *)
  wire _02638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10744" *)
  wire _02639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10744" *)
  wire _02640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10789" *)
  wire _02641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10892" *)
  wire _02642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10921" *)
  wire _02643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11012" *)
  wire _02644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11029" *)
  wire _02645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11138" *)
  wire _02646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11155" *)
  wire _02647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11218" *)
  wire _02648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12028" *)
  wire _02649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12030" *)
  wire _02650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12031" *)
  wire _02651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12031" *)
  wire _02652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12050" *)
  wire _02653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12050" *)
  wire _02654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12052" *)
  wire _02655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12052" *)
  wire _02656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12052" *)
  wire _02657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12053" *)
  wire _02658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12053" *)
  wire _02659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12055" *)
  wire _02660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12056" *)
  wire _02661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12056" *)
  wire _02662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12056" *)
  wire _02663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12060" *)
  wire _02664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12060" *)
  wire _02665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12060" *)
  wire _02666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12078" *)
  wire _02667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12078" *)
  wire _02668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12078" *)
  wire _02669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12098" *)
  wire _02670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12101" *)
  wire _02671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12101" *)
  wire _02672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12108" *)
  wire _02673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12116" *)
  wire _02674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12117" *)
  wire _02675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12117" *)
  wire _02676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12118" *)
  wire _02677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12118" *)
  wire _02678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12120" *)
  wire _02679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12120" *)
  wire _02680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12121" *)
  wire _02681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12121" *)
  wire _02682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12123" *)
  wire _02683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12124" *)
  wire _02684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12124" *)
  wire _02685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12124" *)
  wire _02686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12128" *)
  wire _02687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12128" *)
  wire _02688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12128" *)
  wire _02689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12144" *)
  wire _02690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12157" *)
  wire _02691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12160" *)
  wire _02692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12160" *)
  wire _02693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12179" *)
  wire _02694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12180" *)
  wire _02695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12180" *)
  wire _02696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12180" *)
  wire _02697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12180" *)
  wire _02698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12182" *)
  wire _02699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12182" *)
  wire _02700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12182" *)
  wire _02701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12183" *)
  wire _02702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12183" *)
  wire _02703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12185" *)
  wire _02704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12186" *)
  wire _02705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12186" *)
  wire _02706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12186" *)
  wire _02707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12190" *)
  wire _02708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12190" *)
  wire _02709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12190" *)
  wire _02710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12205" *)
  wire _02711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12208" *)
  wire _02712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12208" *)
  wire _02713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12208" *)
  wire _02714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12222" *)
  wire _02715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12225" *)
  wire _02716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12225" *)
  wire _02717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12244" *)
  wire _02718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12245" *)
  wire _02719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12245" *)
  wire _02720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12246" *)
  wire _02721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12246" *)
  wire _02722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12248" *)
  wire _02723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12248" *)
  wire _02724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12249" *)
  wire _02725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12249" *)
  wire _02726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12251" *)
  wire _02727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12252" *)
  wire _02728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12252" *)
  wire _02729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12252" *)
  wire _02730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12256" *)
  wire _02731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12256" *)
  wire _02732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12256" *)
  wire _02733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12274" *)
  wire _02734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12274" *)
  wire _02735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12281" *)
  wire _02736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12284" *)
  wire _02737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12287" *)
  wire _02738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12288" *)
  wire _02739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12290" *)
  wire _02740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12293" *)
  wire _02741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12302" *)
  wire _02742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12305" *)
  wire _02743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12308" *)
  wire _02744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12309" *)
  wire _02745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12311" *)
  wire _02746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12314" *)
  wire _02747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12323" *)
  wire _02748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12328" *)
  wire _02749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12329" *)
  wire _02750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12331" *)
  wire _02751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12342" *)
  wire _02752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12345" *)
  wire _02753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12348" *)
  wire _02754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12349" *)
  wire _02755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12351" *)
  wire _02756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12354" *)
  wire _02757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12375" *)
  wire _02758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12376" *)
  wire _02759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12376" *)
  wire _02760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12377" *)
  wire _02761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12377" *)
  wire _02762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12377" *)
  wire _02763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12379" *)
  wire _02764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12379" *)
  wire _02765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12380" *)
  wire _02766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12380" *)
  wire _02767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12380" *)
  wire _02768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12383" *)
  wire _02769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12384" *)
  wire _02770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12384" *)
  wire _02771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12384" *)
  wire _02772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12386" *)
  wire _02773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12386" *)
  wire _02774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12386" *)
  wire _02775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12388" *)
  wire _02776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12389" *)
  wire _02777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12389" *)
  wire _02778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12392" *)
  wire _02779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12393" *)
  wire _02780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12393" *)
  wire _02781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12393" *)
  wire _02782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12394" *)
  wire _02783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12401" *)
  wire _02784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12401" *)
  wire _02785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12402" *)
  wire _02786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12402" *)
  wire _02787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12404" *)
  wire _02788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12404" *)
  wire _02789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12405" *)
  wire _02790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12406" *)
  wire _02791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12406" *)
  wire _02792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12409" *)
  wire _02793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12409" *)
  wire _02794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12409" *)
  wire _02795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12411" *)
  wire _02796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12412" *)
  wire _02797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12412" *)
  wire _02798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12414" *)
  wire _02799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12415" *)
  wire _02800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12415" *)
  wire _02801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12422" *)
  wire _02802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12422" *)
  wire _02803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12424" *)
  wire _02804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12424" *)
  wire _02805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12424" *)
  wire _02806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12424" *)
  wire _02807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12426" *)
  wire _02808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12426" *)
  wire _02809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12427" *)
  wire _02810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12427" *)
  wire _02811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12427" *)
  wire _02812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12430" *)
  wire _02813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12430" *)
  wire _02814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12430" *)
  wire _02815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12430" *)
  wire _02816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12432" *)
  wire _02817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12432" *)
  wire _02818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12432" *)
  wire _02819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12435" *)
  wire _02820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12435" *)
  wire _02821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12436" *)
  wire _02822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12436" *)
  wire _02823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12438" *)
  wire _02824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12438" *)
  wire _02825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12438" *)
  wire _02826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12439" *)
  wire _02827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12440" *)
  wire _02828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12440" *)
  wire _02829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12445" *)
  wire _02830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12445" *)
  wire _02831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12448" *)
  wire _02832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12450" *)
  wire _02833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12458" *)
  wire _02834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12458" *)
  wire _02835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12459" *)
  wire _02836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12459" *)
  wire _02837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12461" *)
  wire _02838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12461" *)
  wire _02839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12462" *)
  wire _02840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12462" *)
  wire _02841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12462" *)
  wire _02842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12464" *)
  wire _02843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12467" *)
  wire _02844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12467" *)
  wire _02845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12467" *)
  wire _02846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12477" *)
  wire _02847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12478" *)
  wire _02848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12478" *)
  wire _02849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12479" *)
  wire _02850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12479" *)
  wire _02851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12479" *)
  wire _02852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12481" *)
  wire _02853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12481" *)
  wire _02854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12482" *)
  wire _02855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12482" *)
  wire _02856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12482" *)
  wire _02857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12485" *)
  wire _02858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12486" *)
  wire _02859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12486" *)
  wire _02860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12486" *)
  wire _02861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12488" *)
  wire _02862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12488" *)
  wire _02863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12488" *)
  wire _02864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12490" *)
  wire _02865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12491" *)
  wire _02866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12491" *)
  wire _02867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12494" *)
  wire _02868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12495" *)
  wire _02869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12495" *)
  wire _02870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12495" *)
  wire _02871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12496" *)
  wire _02872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12499" *)
  wire _02873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12499" *)
  wire _02874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12500" *)
  wire _02875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12500" *)
  wire _02876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12502" *)
  wire _02877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12502" *)
  wire _02878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12503" *)
  wire _02879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12504" *)
  wire _02880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12504" *)
  wire _02881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12507" *)
  wire _02882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12507" *)
  wire _02883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12509" *)
  wire _02884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12510" *)
  wire _02885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12512" *)
  wire _02886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12513" *)
  wire _02887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12513" *)
  wire _02888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12520" *)
  wire _02889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12521" *)
  wire _02890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12521" *)
  wire _02891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12522" *)
  wire _02892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12522" *)
  wire _02893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12522" *)
  wire _02894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12524" *)
  wire _02895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12524" *)
  wire _02896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12525" *)
  wire _02897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12525" *)
  wire _02898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12525" *)
  wire _02899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12528" *)
  wire _02900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12529" *)
  wire _02901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12529" *)
  wire _02902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12529" *)
  wire _02903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12531" *)
  wire _02904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12531" *)
  wire _02905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12531" *)
  wire _02906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12533" *)
  wire _02907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12534" *)
  wire _02908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12534" *)
  wire _02909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12537" *)
  wire _02910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12538" *)
  wire _02911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12538" *)
  wire _02912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12538" *)
  wire _02913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12539" *)
  wire _02914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12542" *)
  wire _02915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12542" *)
  wire _02916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12543" *)
  wire _02917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12543" *)
  wire _02918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12545" *)
  wire _02919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12545" *)
  wire _02920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12546" *)
  wire _02921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12546" *)
  wire _02922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12546" *)
  wire _02923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12549" *)
  wire _02924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12549" *)
  wire _02925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12551" *)
  wire _02926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12552" *)
  wire _02927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12554" *)
  wire _02928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12555" *)
  wire _02929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12555" *)
  wire _02930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12560" *)
  wire _02931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12562" *)
  wire _02932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12562" *)
  wire _02933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12566" *)
  wire _02934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12568" *)
  wire _02935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12568" *)
  wire _02936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12572" *)
  wire _02937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12574" *)
  wire _02938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12574" *)
  wire _02939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12578" *)
  wire _02940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12580" *)
  wire _02941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12580" *)
  wire _02942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12622" *)
  wire _02943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12622" *)
  wire _02944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12651" *)
  wire _02945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12692" *)
  wire _02946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12692" *)
  wire _02947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12693" *)
  wire _02948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12695" *)
  wire _02949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12699" *)
  wire _02950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12704" *)
  wire _02951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12706" *)
  wire _02952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12706" *)
  wire _02953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12713" *)
  wire _02954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12713" *)
  wire _02955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12714" *)
  wire _02956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12716" *)
  wire _02957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12722" *)
  wire _02958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12724" *)
  wire _02959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12724" *)
  wire _02960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12730" *)
  wire _02961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12730" *)
  wire _02962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12731" *)
  wire _02963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12733" *)
  wire _02964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12739" *)
  wire _02965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12741" *)
  wire _02966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12741" *)
  wire _02967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12747" *)
  wire _02968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12749" *)
  wire _02969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12754" *)
  wire _02970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12756" *)
  wire _02971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12758" *)
  wire _02972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12758" *)
  wire _02973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12764" *)
  wire _02974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12764" *)
  wire _02975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12765" *)
  wire _02976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12768" *)
  wire _02977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12768" *)
  wire _02978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12769" *)
  wire _02979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12773" *)
  wire _02980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12773" *)
  wire _02981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12781" *)
  wire _02982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12781" *)
  wire _02983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12782" *)
  wire _02984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12801" *)
  wire _02985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12801" *)
  wire _02986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12804" *)
  wire _02987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12804" *)
  wire _02988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12807" *)
  wire _02989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12807" *)
  wire _02990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12808" *)
  wire _02991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12808" *)
  wire _02992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12809" *)
  wire _02993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12809" *)
  wire _02994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12811" *)
  wire _02995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12812" *)
  wire _02996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12812" *)
  wire _02997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12813" *)
  wire _02998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12813" *)
  wire _02999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12814" *)
  wire _03000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12815" *)
  wire _03001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12824" *)
  wire _03002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12833" *)
  wire _03003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12835" *)
  wire _03004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12836" *)
  wire _03005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12837" *)
  wire _03006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12860" *)
  wire _03007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12860" *)
  wire _03008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12861" *)
  wire _03009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12861" *)
  wire _03010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12862" *)
  wire _03011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12864" *)
  wire _03012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12864" *)
  wire _03013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12865" *)
  wire _03014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12865" *)
  wire _03015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *)
  wire _03016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12873" *)
  wire _03017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12880" *)
  wire _03018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12883" *)
  wire _03019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12883" *)
  wire _03020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12907" *)
  wire _03021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12907" *)
  wire _03022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12908" *)
  wire _03023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12908" *)
  wire _03024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12909" *)
  wire _03025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12909" *)
  wire _03026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12911" *)
  wire _03027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12911" *)
  wire _03028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12912" *)
  wire _03029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12912" *)
  wire _03030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *)
  wire _03031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12920" *)
  wire _03032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12927" *)
  wire _03033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12929" *)
  wire _03034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12930" *)
  wire _03035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12930" *)
  wire _03036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12932" *)
  wire _03037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12932" *)
  wire _03038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12939" *)
  wire _03039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12944" *)
  wire _03040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12944" *)
  wire _03041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12945" *)
  wire _03042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12967" *)
  wire _03043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12967" *)
  wire _03044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12968" *)
  wire _03045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12968" *)
  wire _03046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12969" *)
  wire _03047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12969" *)
  wire _03048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12971" *)
  wire _03049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12971" *)
  wire _03050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12972" *)
  wire _03051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12972" *)
  wire _03052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12973" *)
  wire _03053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12973" *)
  wire _03054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12974" *)
  wire _03055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12988" *)
  wire _03056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12990" *)
  wire _03057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12991" *)
  wire _03058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12991" *)
  wire _03059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12993" *)
  wire _03060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12993" *)
  wire _03061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12998" *)
  wire _03062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12998" *)
  wire _03063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12999" *)
  wire _03064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13000" *)
  wire _03065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13001" *)
  wire _03066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13001" *)
  wire _03067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13005" *)
  wire _03068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13005" *)
  wire _03069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13015" *)
  wire _03070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13016" *)
  wire _03071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13018" *)
  wire _03072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13018" *)
  wire _03073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13022" *)
  wire _03074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13022" *)
  wire _03075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13031" *)
  wire _03076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13032" *)
  wire _03077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13034" *)
  wire _03078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13034" *)
  wire _03079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13038" *)
  wire _03080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13038" *)
  wire _03081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13047" *)
  wire _03082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13048" *)
  wire _03083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13050" *)
  wire _03084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13050" *)
  wire _03085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13054" *)
  wire _03086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13054" *)
  wire _03087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13064" *)
  wire _03088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13065" *)
  wire _03089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13065" *)
  wire _03090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13067" *)
  wire _03091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13067" *)
  wire _03092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13067" *)
  wire _03093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13069" *)
  wire _03094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13069" *)
  wire _03095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13070" *)
  wire _03096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13070" *)
  wire _03097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13073" *)
  wire _03098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13074" *)
  wire _03099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13076" *)
  wire _03100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13079" *)
  wire _03101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13079" *)
  wire _03102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13081" *)
  wire _03103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13081" *)
  wire _03104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13083" *)
  wire _03105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13084" *)
  wire _03106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13084" *)
  wire _03107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13086" *)
  wire _03108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13086" *)
  wire _03109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13088" *)
  wire _03110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13090" *)
  wire _03111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13090" *)
  wire _03112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13090" *)
  wire _03113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13092" *)
  wire _03114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13093" *)
  wire _03115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13093" *)
  wire _03116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13095" *)
  wire _03117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13095" *)
  wire _03118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13097" *)
  wire _03119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13099" *)
  wire _03120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13099" *)
  wire _03121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13101" *)
  wire _03122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13102" *)
  wire _03123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13102" *)
  wire _03124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13104" *)
  wire _03125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13104" *)
  wire _03126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13106" *)
  wire _03127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13107" *)
  wire _03128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13107" *)
  wire _03129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13109" *)
  wire _03130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13111" *)
  wire _03131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13111" *)
  wire _03132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13112" *)
  wire _03133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13112" *)
  wire _03134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13116" *)
  wire _03135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13118" *)
  wire _03136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13118" *)
  wire _03137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13118" *)
  wire _03138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13121" *)
  wire _03139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13121" *)
  wire _03140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13123" *)
  wire _03141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13123" *)
  wire _03142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13125" *)
  wire _03143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13126" *)
  wire _03144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13126" *)
  wire _03145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13128" *)
  wire _03146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13128" *)
  wire _03147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13134" *)
  wire _03148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13134" *)
  wire _03149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13139" *)
  wire _03150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13139" *)
  wire _03151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13139" *)
  wire _03152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13147" *)
  wire _03153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13153" *)
  wire _03154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13170" *)
  wire _03155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13180" *)
  wire _03156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13186" *)
  wire _03157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13186" *)
  wire _03158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13190" *)
  wire _03159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13190" *)
  wire _03160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13190" *)
  wire _03161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13209" *)
  wire _03162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13214" *)
  wire _03163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13214" *)
  wire _03164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13214" *)
  wire _03165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13219" *)
  wire _03166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13219" *)
  wire _03167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13219" *)
  wire _03168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13221" *)
  wire _03169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13236" *)
  wire _03170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13249" *)
  wire _03171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13262" *)
  wire _03172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13273" *)
  wire _03173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13273" *)
  wire _03174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *)
  wire _03188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *)
  wire _03202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _03203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _03204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _03205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _03206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _03207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _03208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _03209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *)
  wire _03210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _03211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _03212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _03213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _03214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _03215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _03216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _03217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *)
  wire _03218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _03219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _03220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _03221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _03222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _03223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _03224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _03225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *)
  wire _03226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *)
  wire [11:0] _03227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *)
  wire [11:0] _03228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *)
  wire [11:0] _03229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *)
  wire [11:0] _03230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *)
  wire [11:0] _03231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *)
  wire [11:0] _03232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *)
  wire [11:0] _03233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *)
  wire [11:0] _03234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *)
  wire [11:0] _03235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *)
  wire [11:0] _03236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *)
  wire [11:0] _03237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *)
  wire [11:0] _03238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *)
  wire [22:0] _03239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *)
  wire [22:0] _03240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *)
  wire [22:0] _03241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *)
  wire [22:0] _03242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *)
  wire [22:0] _03243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *)
  wire [22:0] _03244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *)
  wire [22:0] _03245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *)
  wire [22:0] _03246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *)
  wire [22:0] _03247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *)
  wire [22:0] _03248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *)
  wire [22:0] _03249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *)
  wire [22:0] _03250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *)
  wire [22:0] _03251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *)
  wire [22:0] _03252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *)
  wire [22:0] _03253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *)
  wire [22:0] _03254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *)
  wire [22:0] _03255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *)
  wire [22:0] _03256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *)
  wire [22:0] _03257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *)
  wire [22:0] _03258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *)
  wire [1:0] _03259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *)
  wire [1:0] _03260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *)
  wire [1:0] _03261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *)
  wire [1:0] _03262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *)
  wire [1:0] _03263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *)
  wire [1:0] _03264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *)
  wire [1:0] _03265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *)
  wire [1:0] _03266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *)
  wire [49:0] _03267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *)
  wire [49:0] _03268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *)
  wire [49:0] _03269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *)
  wire [49:0] _03270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *)
  wire [49:0] _03271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *)
  wire [49:0] _03272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *)
  wire [49:0] _03273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *)
  wire [49:0] _03274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *)
  wire [49:0] _03275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *)
  wire [49:0] _03276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *)
  wire [49:0] _03277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *)
  wire [49:0] _03278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *)
  wire [5:0] _03279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *)
  wire [5:0] _03280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *)
  wire [5:0] _03281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *)
  wire [5:0] _03282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *)
  wire [5:0] _03283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *)
  wire [5:0] _03284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *)
  wire [5:0] _03285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *)
  wire [5:0] _03286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *)
  wire [5:0] _03287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *)
  wire [5:0] _03288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *)
  wire [5:0] _03289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *)
  wire [5:0] _03290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *)
  wire [5:0] _03291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *)
  wire [5:0] _03292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *)
  wire [5:0] _03293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *)
  wire [5:0] _03294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *)
  wire [5:0] _03295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *)
  wire [5:0] _03296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *)
  wire [5:0] _03297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *)
  wire [5:0] _03298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *)
  wire [5:0] _03299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *)
  wire [5:0] _03300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *)
  wire [5:0] _03301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *)
  wire [5:0] _03302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *)
  wire [5:0] _03303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *)
  wire [5:0] _03304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *)
  wire [5:0] _03305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *)
  wire [5:0] _03306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *)
  wire [7:0] _03307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *)
  wire [7:0] _03308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *)
  wire [7:0] _03309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *)
  wire [7:0] _03310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *)
  wire [7:0] _03311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *)
  wire [7:0] _03312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *)
  wire [7:0] _03313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *)
  wire [7:0] _03314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _03315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _03316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _03317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _03318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _03319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _03320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _03321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *)
  wire [7:0] _03322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _03323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _03324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _03325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _03326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _03327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _03328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _03329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *)
  wire [7:0] _03330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _03331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _03332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _03333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _03334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _03335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _03336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _03337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *)
  wire [7:0] _03338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *)
  wire [8:0] _03339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *)
  wire [8:0] _03340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *)
  wire [8:0] _03341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *)
  wire [8:0] _03342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13446" *)
  wire [8:0] _03343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13446" *)
  wire [8:0] _03344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13446" *)
  wire [8:0] _03345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13446" *)
  wire [8:0] _03346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *)
  wire [8:0] _03347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *)
  wire [8:0] _03348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *)
  wire [8:0] _03349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *)
  wire [8:0] _03350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5452" *)
  wire _03351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5454" *)
  wire _03352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5456" *)
  wire _03353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5458" *)
  wire _03354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5460" *)
  wire _03355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5475" *)
  wire _03356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5496" *)
  wire _03357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5503" *)
  wire _03358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5512" *)
  wire _03359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5532" *)
  wire _03360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5533" *)
  wire _03361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5533" *)
  wire _03362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5533" *)
  wire _03363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5533" *)
  wire _03364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5535" *)
  wire _03365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5535" *)
  wire _03366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5535" *)
  wire _03367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5536" *)
  wire _03368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5536" *)
  wire _03369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5540" *)
  wire _03370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5556" *)
  wire _03371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5556" *)
  wire _03372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5558" *)
  wire _03373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5564" *)
  wire _03374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5568" *)
  wire _03375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5579" *)
  wire _03376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5580" *)
  wire _03377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5581" *)
  wire _03378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5581" *)
  wire _03379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5582" *)
  wire _03380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5582" *)
  wire _03381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5584" *)
  wire _03382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5584" *)
  wire _03383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5585" *)
  wire _03384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5585" *)
  wire _03385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5590" *)
  wire _03386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5606" *)
  wire _03387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5606" *)
  wire _03388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5611" *)
  wire _03389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5613" *)
  wire _03390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5621" *)
  wire _03391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5622" *)
  wire _03392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5622" *)
  wire _03393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5623" *)
  wire _03394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5623" *)
  wire _03395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5625" *)
  wire _03396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5625" *)
  wire _03397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5626" *)
  wire _03398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5626" *)
  wire _03399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5630" *)
  wire _03400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5644" *)
  wire _03401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5647" *)
  wire _03402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5652" *)
  wire _03403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5653" *)
  wire _03404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5653" *)
  wire _03405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5654" *)
  wire _03406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5654" *)
  wire _03407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5656" *)
  wire _03408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5656" *)
  wire _03409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5657" *)
  wire _03410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5657" *)
  wire _03411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5661" *)
  wire _03412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5675" *)
  wire _03413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5677" *)
  wire _03414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5687" *)
  wire _03415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5688" *)
  wire _03416_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5692" *)
  wire _03417_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5693" *)
  wire _03418_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5693" *)
  wire _03419_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5693" *)
  wire _03420_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5693" *)
  wire _03421_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5695" *)
  wire _03422_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5695" *)
  wire _03423_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5695" *)
  wire _03424_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5702" *)
  wire _03425_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5707" *)
  wire _03426_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5707" *)
  wire _03427_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5707" *)
  wire _03428_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5708" *)
  wire _03429_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5708" *)
  wire _03430_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5710" *)
  wire _03431_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5710" *)
  wire _03432_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5720" *)
  wire _03433_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5720" *)
  wire _03434_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5720" *)
  wire _03435_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5721" *)
  wire _03436_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5721" *)
  wire _03437_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5723" *)
  wire _03438_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5723" *)
  wire _03439_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5723" *)
  wire _03440_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5731" *)
  wire _03441_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5731" *)
  wire _03442_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5732" *)
  wire _03443_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5732" *)
  wire _03444_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5732" *)
  wire _03445_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5734" *)
  wire _03446_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5734" *)
  wire _03447_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5734" *)
  wire _03448_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5776" *)
  wire _03449_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5780" *)
  wire _03450_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5786" *)
  wire _03451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5814" *)
  wire _03452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5814" *)
  wire _03453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5821" *)
  wire _03454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5841" *)
  wire _03455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5845" *)
  wire _03456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5846" *)
  wire _03457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5905" *)
  wire _03458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5905" *)
  wire _03459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5912" *)
  wire _03460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5926" *)
  wire _03461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5944" *)
  wire _03462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5964" *)
  wire _03463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5965" *)
  wire _03464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5966" *)
  wire _03465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5975" *)
  wire _03466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5975" *)
  wire _03467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5977" *)
  wire _03468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5977" *)
  wire _03469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5980" *)
  wire _03470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5982" *)
  wire _03471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6013" *)
  wire _03472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6013" *)
  wire _03473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6014" *)
  wire _03474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6033" *)
  wire _03475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6033" *)
  wire _03476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6035" *)
  wire _03477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6035" *)
  wire _03478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6038" *)
  wire _03479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6040" *)
  wire _03480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6059" *)
  wire _03481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6059" *)
  wire _03482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6060" *)
  wire _03483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6078" *)
  wire _03484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6078" *)
  wire _03485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6080" *)
  wire _03486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6080" *)
  wire _03487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6083" *)
  wire _03488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6085" *)
  wire _03489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6085" *)
  wire _03490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6120" *)
  wire _03491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6120" *)
  wire _03492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6121" *)
  wire _03493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6124" *)
  wire _03494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6125" *)
  wire _03495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6131" *)
  wire _03496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6158" *)
  wire _03497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6158" *)
  wire _03498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6160" *)
  wire _03499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6160" *)
  wire _03500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6166" *)
  wire _03501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6168" *)
  wire _03502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6191" *)
  wire _03503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6192" *)
  wire _03504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6199" *)
  wire _03505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6199" *)
  wire _03506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6200" *)
  wire _03507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6200" *)
  wire _03508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6201" *)
  wire _03509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6201" *)
  wire _03510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6202" *)
  wire _03511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6202" *)
  wire _03512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6203" *)
  wire _03513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6203" *)
  wire _03514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6204" *)
  wire _03515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6204" *)
  wire _03516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6205" *)
  wire _03517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6205" *)
  wire _03518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6206" *)
  wire _03519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6206" *)
  wire _03520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6207" *)
  wire _03521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6207" *)
  wire _03522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6208" *)
  wire _03523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6208" *)
  wire _03524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6209" *)
  wire _03525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6209" *)
  wire _03526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6210" *)
  wire _03527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6210" *)
  wire _03528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6219" *)
  wire _03529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6219" *)
  wire _03530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6220" *)
  wire _03531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6220" *)
  wire _03532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6221" *)
  wire _03533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6221" *)
  wire _03534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6222" *)
  wire _03535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6222" *)
  wire _03536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6223" *)
  wire _03537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6223" *)
  wire _03538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6224" *)
  wire _03539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6224" *)
  wire _03540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6225" *)
  wire _03541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6225" *)
  wire _03542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6226" *)
  wire _03543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6226" *)
  wire _03544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6227" *)
  wire _03545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6227" *)
  wire _03546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6228" *)
  wire _03547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6228" *)
  wire _03548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6229" *)
  wire _03549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6229" *)
  wire _03550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6230" *)
  wire _03551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6230" *)
  wire _03552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6239" *)
  wire _03553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6239" *)
  wire _03554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6240" *)
  wire _03555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6240" *)
  wire _03556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6241" *)
  wire _03557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6241" *)
  wire _03558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6242" *)
  wire _03559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6242" *)
  wire _03560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6243" *)
  wire _03561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6243" *)
  wire _03562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6244" *)
  wire _03563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6244" *)
  wire _03564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6245" *)
  wire _03565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6245" *)
  wire _03566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6246" *)
  wire _03567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6246" *)
  wire _03568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6247" *)
  wire _03569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6247" *)
  wire _03570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6248" *)
  wire _03571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6248" *)
  wire _03572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6249" *)
  wire _03573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6249" *)
  wire _03574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6250" *)
  wire _03575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6250" *)
  wire _03576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6259" *)
  wire _03577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6259" *)
  wire _03578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6260" *)
  wire _03579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6260" *)
  wire _03580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6261" *)
  wire _03581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6261" *)
  wire _03582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6262" *)
  wire _03583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6262" *)
  wire _03584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6263" *)
  wire _03585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6263" *)
  wire _03586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6264" *)
  wire _03587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6264" *)
  wire _03588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6265" *)
  wire _03589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6265" *)
  wire _03590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6266" *)
  wire _03591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6266" *)
  wire _03592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6267" *)
  wire _03593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6267" *)
  wire _03594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6268" *)
  wire _03595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6268" *)
  wire _03596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6269" *)
  wire _03597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6269" *)
  wire _03598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6270" *)
  wire _03599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6270" *)
  wire _03600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6279" *)
  wire _03601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6279" *)
  wire _03602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6280" *)
  wire _03603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6280" *)
  wire _03604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6281" *)
  wire _03605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6281" *)
  wire _03606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6282" *)
  wire _03607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6282" *)
  wire _03608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6283" *)
  wire _03609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6283" *)
  wire _03610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6284" *)
  wire _03611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6284" *)
  wire _03612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6285" *)
  wire _03613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6285" *)
  wire _03614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6286" *)
  wire _03615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6286" *)
  wire _03616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6287" *)
  wire _03617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6287" *)
  wire _03618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6288" *)
  wire _03619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6288" *)
  wire _03620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6289" *)
  wire _03621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6289" *)
  wire _03622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6290" *)
  wire _03623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6290" *)
  wire _03624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6299" *)
  wire _03625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6299" *)
  wire _03626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6300" *)
  wire _03627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6300" *)
  wire _03628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6301" *)
  wire _03629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6301" *)
  wire _03630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6302" *)
  wire _03631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6302" *)
  wire _03632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6303" *)
  wire _03633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6303" *)
  wire _03634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6304" *)
  wire _03635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6304" *)
  wire _03636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6305" *)
  wire _03637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6305" *)
  wire _03638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6306" *)
  wire _03639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6306" *)
  wire _03640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6307" *)
  wire _03641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6307" *)
  wire _03642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6308" *)
  wire _03643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6308" *)
  wire _03644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6309" *)
  wire _03645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6309" *)
  wire _03646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6310" *)
  wire _03647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6310" *)
  wire _03648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6319" *)
  wire _03649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6319" *)
  wire _03650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6320" *)
  wire _03651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6320" *)
  wire _03652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6321" *)
  wire _03653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6321" *)
  wire _03654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6322" *)
  wire _03655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6322" *)
  wire _03656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6323" *)
  wire _03657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6323" *)
  wire _03658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6324" *)
  wire _03659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6324" *)
  wire _03660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6325" *)
  wire _03661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6325" *)
  wire _03662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6326" *)
  wire _03663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6326" *)
  wire _03664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6327" *)
  wire _03665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6327" *)
  wire _03666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6328" *)
  wire _03667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6328" *)
  wire _03668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6329" *)
  wire _03669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6329" *)
  wire _03670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6330" *)
  wire _03671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6330" *)
  wire _03672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6339" *)
  wire _03673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6339" *)
  wire _03674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6340" *)
  wire _03675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6340" *)
  wire _03676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6341" *)
  wire _03677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6341" *)
  wire _03678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6342" *)
  wire _03679_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6342" *)
  wire _03680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6343" *)
  wire _03681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6343" *)
  wire _03682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6344" *)
  wire _03683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6344" *)
  wire _03684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6345" *)
  wire _03685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6345" *)
  wire _03686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6346" *)
  wire _03687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6346" *)
  wire _03688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6347" *)
  wire _03689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6347" *)
  wire _03690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6348" *)
  wire _03691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6348" *)
  wire _03692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6349" *)
  wire _03693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6349" *)
  wire _03694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6350" *)
  wire _03695_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6350" *)
  wire _03696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6358" *)
  wire _03697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6368" *)
  wire _03698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6374" *)
  wire _03699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6381" *)
  wire _03700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6389" *)
  wire _03701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6396" *)
  wire _03702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6404" *)
  wire _03703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6411" *)
  wire _03704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6477" *)
  wire _03705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6478" *)
  wire _03706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6483" *)
  wire _03707_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6484" *)
  wire _03708_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6486" *)
  wire _03709_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6487" *)
  wire _03710_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6489" *)
  wire _03711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6549" *)
  wire _03712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6595" *)
  wire _03713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6609" *)
  wire _03714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6623" *)
  wire _03715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6646" *)
  wire _03716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6660" *)
  wire _03717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6676" *)
  wire _03718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6699" *)
  wire _03719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6713" *)
  wire _03720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6727" *)
  wire _03721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6750" *)
  wire _03722_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6764" *)
  wire _03723_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6778" *)
  wire _03724_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6867" *)
  wire _03725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6925" *)
  wire _03726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6983" *)
  wire _03727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7041" *)
  wire _03728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7073" *)
  wire _03729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7081" *)
  wire _03730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7083" *)
  wire _03731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7084" *)
  wire _03732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7085" *)
  wire _03733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7095" *)
  wire _03734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7097" *)
  wire _03735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7098" *)
  wire _03736_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7099" *)
  wire _03737_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7109" *)
  wire _03738_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7111" *)
  wire _03739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7112" *)
  wire _03740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7113" *)
  wire _03741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7123" *)
  wire _03742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7125" *)
  wire _03743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7126" *)
  wire _03744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7127" *)
  wire _03745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7456" *)
  wire _03746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7458" *)
  wire _03747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7460" *)
  wire _03748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7462" *)
  wire _03749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7464" *)
  wire _03750_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7472" *)
  wire _03751_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7472" *)
  wire _03752_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7484" *)
  wire _03753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7490" *)
  wire _03754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7498" *)
  wire _03755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7511" *)
  wire _03756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7511" *)
  wire _03757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7524" *)
  wire _03758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7524" *)
  wire _03759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7524" *)
  wire _03760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7532" *)
  wire _03761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7536" *)
  wire _03762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7537" *)
  wire _03763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7537" *)
  wire _03764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7543" *)
  wire _03765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7544" *)
  wire _03766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7548" *)
  wire _03767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7549" *)
  wire _03768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7551" *)
  wire _03769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7553" *)
  wire _03770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7553" *)
  wire _03771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7557" *)
  wire _03772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7557" *)
  wire _03773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7566" *)
  wire _03774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7567" *)
  wire _03775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7569" *)
  wire _03776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7569" *)
  wire _03777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7572" *)
  wire _03778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7572" *)
  wire _03779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7575" *)
  wire _03780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7575" *)
  wire _03781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7577" *)
  wire _03782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7577" *)
  wire _03783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7580" *)
  wire _03784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7580" *)
  wire _03785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7581" *)
  wire _03786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7584" *)
  wire _03787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7586" *)
  wire _03788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7587" *)
  wire _03789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7595" *)
  wire _03790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7595" *)
  wire _03791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7604" *)
  wire _03792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7613" *)
  wire _03793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7616" *)
  wire _03794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7620" *)
  wire _03795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7622" *)
  wire _03796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7623" *)
  wire _03797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7633" *)
  wire _03798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *)
  wire _03799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *)
  wire _03800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *)
  wire _03801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7651" *)
  wire _03802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7651" *)
  wire _03803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7661" *)
  wire _03804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7665" *)
  wire _03805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7669" *)
  wire _03806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7690" *)
  wire _03807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7690" *)
  wire _03808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7697" *)
  wire _03809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7697" *)
  wire _03810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7705" *)
  wire _03811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7705" *)
  wire _03812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7713" *)
  wire _03813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7713" *)
  wire _03814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7723" *)
  wire _03815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7725" *)
  wire _03816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7727" *)
  wire _03817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7729" *)
  wire _03818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7731" *)
  wire _03819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7733" *)
  wire _03820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7735" *)
  wire _03821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7737" *)
  wire _03822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7754" *)
  wire _03823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7759" *)
  wire _03824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7764" *)
  wire _03825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7769" *)
  wire _03826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7814" *)
  wire _03827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7817" *)
  wire _03828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7822" *)
  wire _03829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7823" *)
  wire _03830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7823" *)
  wire _03831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7827" *)
  wire _03832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7831" *)
  wire _03833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7836" *)
  wire _03834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7838" *)
  wire _03835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7843" *)
  wire _03836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7847" *)
  wire _03837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7848" *)
  wire _03838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7849" *)
  wire _03839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7851" *)
  wire _03840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7852" *)
  wire _03841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7852" *)
  wire _03842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7856" *)
  wire _03843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7856" *)
  wire _03844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7856" *)
  wire _03845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7860" *)
  wire _03846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7861" *)
  wire _03847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7861" *)
  wire _03848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7864" *)
  wire _03849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7869" *)
  wire _03850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7869" *)
  wire _03851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8086" *)
  wire _03852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8094" *)
  wire _03853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8197" *)
  wire _03854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8211" *)
  wire _03855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8217" *)
  wire _03856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8224" *)
  wire _03857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8278" *)
  wire _03858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8286" *)
  wire _03859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8286" *)
  wire _03860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8286" *)
  wire _03861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8311" *)
  wire _03862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8333" *)
  wire _03863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8341" *)
  wire _03864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8341" *)
  wire _03865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8341" *)
  wire _03866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8364" *)
  wire _03867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8373" *)
  wire _03868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8382" *)
  wire _03869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8382" *)
  wire _03870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8382" *)
  wire _03871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8413" *)
  wire _03872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8422" *)
  wire _03873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8431" *)
  wire _03874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8431" *)
  wire _03875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8431" *)
  wire _03876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8444" *)
  wire _03877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8453" *)
  wire _03878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8503" *)
  wire _03879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8503" *)
  wire _03880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8526" *)
  wire _03881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8676" *)
  wire _03882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8676" *)
  wire _03883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8746" *)
  wire _03884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8835" *)
  wire _03885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8835" *)
  wire _03886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8894" *)
  wire _03887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8915" *)
  wire _03888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8915" *)
  wire _03889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8916" *)
  wire _03890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8969" *)
  wire _03891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8969" *)
  wire _03892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9014" *)
  wire _03893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9035" *)
  wire _03894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9035" *)
  wire _03895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9036" *)
  wire _03896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9089" *)
  wire _03897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9089" *)
  wire _03898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9111" *)
  wire _03899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9433" *)
  wire _03900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9589" *)
  wire _03901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9719" *)
  wire _03902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9813" *)
  wire _03903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9911" *)
  wire _03904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5989" *)
  wire _03905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8141" *)
  wire _03906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8155" *)
  wire _03907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8192" *)
  wire _03908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8194" *)
  wire _03909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8196" *)
  wire _03910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8199" *)
  wire _03911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8202" *)
  wire _03912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8204" *)
  wire _03913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1760" *)
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1772" *)
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1768" *)
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1764" *)
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2449" *)
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2444" *)
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2294" *)
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2310" *)
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2326" *)
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2342" *)
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1408" *)
  reg [7:0] FpAdd_8U_23U_1_a_right_shift_qr_1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1376" *)
  reg [7:0] FpAdd_8U_23U_1_a_right_shift_qr_2_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1344" *)
  reg [7:0] FpAdd_8U_23U_1_a_right_shift_qr_3_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1312" *)
  reg [7:0] FpAdd_8U_23U_1_a_right_shift_qr_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2307" *)
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2291" *)
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2339" *)
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2323" *)
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2292" *)
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2308" *)
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2324" *)
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2340" *)
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2293" *)
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2309" *)
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2325" *)
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2341" *)
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1809" *)
  wire FpAdd_8U_23U_1_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1808" *)
  wire FpAdd_8U_23U_1_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3932" *)
  wire FpAdd_8U_23U_1_and_35_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3948" *)
  wire FpAdd_8U_23U_1_and_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3964" *)
  wire FpAdd_8U_23U_1_and_39_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1807" *)
  wire FpAdd_8U_23U_1_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3980" *)
  wire FpAdd_8U_23U_1_and_41_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2535" *)
  wire FpAdd_8U_23U_1_and_46_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2232" *)
  wire FpAdd_8U_23U_1_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1407" *)
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1375" *)
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_2_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1343" *)
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_3_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1311" *)
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2502" *)
  wire FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2503" *)
  wire FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2501" *)
  wire FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1901" *)
  wire FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2651" *)
  wire FpAdd_8U_23U_1_is_a_greater_acc_10_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4089" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpAdd_8U_23U_1_is_a_greater_acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2648" *)
  wire FpAdd_8U_23U_1_is_a_greater_acc_4_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4083" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpAdd_8U_23U_1_is_a_greater_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2649" *)
  wire FpAdd_8U_23U_1_is_a_greater_acc_6_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4085" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpAdd_8U_23U_1_is_a_greater_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2650" *)
  wire FpAdd_8U_23U_1_is_a_greater_acc_8_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4087" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpAdd_8U_23U_1_is_a_greater_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1450" *)
  reg FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1481" *)
  reg FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1511" *)
  reg FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1541" *)
  reg FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2524" *)
  wire FpAdd_8U_23U_1_is_a_greater_oelse_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2474" *)
  wire FpAdd_8U_23U_1_is_addition_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1452" *)
  reg FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1483" *)
  reg FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1513" *)
  reg FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2576" *)
  wire FpAdd_8U_23U_1_is_inf_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1543" *)
  reg FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2563" *)
  wire FpAdd_8U_23U_1_lut_lookup_else_else_else_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2052" *)
  wire [7:0] FpAdd_8U_23U_1_mux1h_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2055" *)
  wire [7:0] FpAdd_8U_23U_1_mux1h_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2058" *)
  wire [7:0] FpAdd_8U_23U_1_mux1h_5_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2061" *)
  wire [7:0] FpAdd_8U_23U_1_mux1h_7_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1579" *)
  reg FpAdd_8U_23U_1_mux_13_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1580" *)
  reg FpAdd_8U_23U_1_mux_13_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1604" *)
  reg FpAdd_8U_23U_1_mux_17_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1578" *)
  reg FpAdd_8U_23U_1_mux_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1605" *)
  reg FpAdd_8U_23U_1_mux_29_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1606" *)
  reg FpAdd_8U_23U_1_mux_29_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1630" *)
  reg FpAdd_8U_23U_1_mux_33_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1631" *)
  reg FpAdd_8U_23U_1_mux_45_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1632" *)
  reg FpAdd_8U_23U_1_mux_45_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1660" *)
  reg FpAdd_8U_23U_1_mux_49_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1661" *)
  reg FpAdd_8U_23U_1_mux_61_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1662" *)
  reg FpAdd_8U_23U_1_mux_61_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1451" *)
  reg [7:0] FpAdd_8U_23U_1_qr_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1482" *)
  reg [7:0] FpAdd_8U_23U_1_qr_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1512" *)
  reg [7:0] FpAdd_8U_23U_1_qr_4_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1542" *)
  reg [7:0] FpAdd_8U_23U_1_qr_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2050" *)
  wire [7:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_11_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2042" *)
  wire [7:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2045" *)
  wire [7:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_5_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2048" *)
  wire [7:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_8_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1758" *)
  wire FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_11_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1770" *)
  wire FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_5_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1766" *)
  wire FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_7_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1762" *)
  wire FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_9_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3890" *)
  wire [22:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3896" *)
  wire [22:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3902" *)
  wire [22:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3908" *)
  wire [22:0] FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2298" *)
  wire [48:0] FpAdd_8U_23U_2_a_int_mant_p1_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2314" *)
  wire [48:0] FpAdd_8U_23U_2_a_int_mant_p1_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2330" *)
  wire [48:0] FpAdd_8U_23U_2_a_int_mant_p1_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2346" *)
  wire [48:0] FpAdd_8U_23U_2_a_int_mant_p1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3271" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3272" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3287" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3288" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3279" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3280" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3295" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3296" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qelse_mux_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2300" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qr_1_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1396" *)
  reg [7:0] FpAdd_8U_23U_2_a_right_shift_qr_1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2316" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qr_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1364" *)
  reg [7:0] FpAdd_8U_23U_2_a_right_shift_qr_2_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2332" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qr_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1332" *)
  reg [7:0] FpAdd_8U_23U_2_a_right_shift_qr_3_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2348" *)
  wire [7:0] FpAdd_8U_23U_2_a_right_shift_qr_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1300" *)
  reg [7:0] FpAdd_8U_23U_2_a_right_shift_qr_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2311" *)
  wire [48:0] FpAdd_8U_23U_2_addend_larger_asn_13_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2295" *)
  wire [48:0] FpAdd_8U_23U_2_addend_larger_asn_19_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2343" *)
  wire [48:0] FpAdd_8U_23U_2_addend_larger_asn_1_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2327" *)
  wire [48:0] FpAdd_8U_23U_2_addend_larger_asn_7_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2296" *)
  wire [48:0] FpAdd_8U_23U_2_addend_larger_qr_1_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2312" *)
  wire [48:0] FpAdd_8U_23U_2_addend_larger_qr_2_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2328" *)
  wire [48:0] FpAdd_8U_23U_2_addend_larger_qr_3_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2344" *)
  wire [48:0] FpAdd_8U_23U_2_addend_larger_qr_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2297" *)
  wire [48:0] FpAdd_8U_23U_2_addend_smaller_qr_1_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2313" *)
  wire [48:0] FpAdd_8U_23U_2_addend_smaller_qr_2_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2329" *)
  wire [48:0] FpAdd_8U_23U_2_addend_smaller_qr_3_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2345" *)
  wire [48:0] FpAdd_8U_23U_2_addend_smaller_qr_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1992" *)
  wire FpAdd_8U_23U_2_and_10_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1993" *)
  wire FpAdd_8U_23U_2_and_11_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3956" *)
  wire FpAdd_8U_23U_2_and_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3958" *)
  wire FpAdd_8U_23U_2_and_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1997" *)
  wire FpAdd_8U_23U_2_and_16_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1998" *)
  wire FpAdd_8U_23U_2_and_17_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3972" *)
  wire FpAdd_8U_23U_2_and_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2236" *)
  wire FpAdd_8U_23U_2_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3974" *)
  wire FpAdd_8U_23U_2_and_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2003" *)
  wire FpAdd_8U_23U_2_and_22_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2004" *)
  wire FpAdd_8U_23U_2_and_23_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3988" *)
  wire FpAdd_8U_23U_2_and_25_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3990" *)
  wire FpAdd_8U_23U_2_and_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3941" *)
  wire FpAdd_8U_23U_2_and_28_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3955" *)
  wire FpAdd_8U_23U_2_and_29_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2238" *)
  wire FpAdd_8U_23U_2_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3957" *)
  wire FpAdd_8U_23U_2_and_30_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3971" *)
  wire FpAdd_8U_23U_2_and_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3973" *)
  wire FpAdd_8U_23U_2_and_32_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3987" *)
  wire FpAdd_8U_23U_2_and_33_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3989" *)
  wire FpAdd_8U_23U_2_and_34_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2436" *)
  wire FpAdd_8U_23U_2_and_35_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2437" *)
  wire FpAdd_8U_23U_2_and_36_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2439" *)
  wire FpAdd_8U_23U_2_and_37_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2240" *)
  wire FpAdd_8U_23U_2_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2518" *)
  wire FpAdd_8U_23U_2_and_44_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1986" *)
  wire FpAdd_8U_23U_2_and_4_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1987" *)
  wire FpAdd_8U_23U_2_and_5_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3940" *)
  wire FpAdd_8U_23U_2_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3942" *)
  wire FpAdd_8U_23U_2_and_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3939" *)
  wire FpAdd_8U_23U_2_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2234" *)
  wire FpAdd_8U_23U_2_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2229" *)
  wire [22:0] FpAdd_8U_23U_2_asn_35_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2228" *)
  wire [22:0] FpAdd_8U_23U_2_asn_40_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2227" *)
  wire [22:0] FpAdd_8U_23U_2_asn_45_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2226" *)
  wire [22:0] FpAdd_8U_23U_2_asn_50_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2170" *)
  wire FpAdd_8U_23U_2_b_right_shift_qif_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2171" *)
  wire FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2174" *)
  wire FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2175" *)
  wire FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2299" *)
  wire [7:0] FpAdd_8U_23U_2_b_right_shift_qr_1_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2315" *)
  wire [7:0] FpAdd_8U_23U_2_b_right_shift_qr_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2331" *)
  wire [7:0] FpAdd_8U_23U_2_b_right_shift_qr_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2347" *)
  wire [7:0] FpAdd_8U_23U_2_b_right_shift_qr_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3936" *)
  wire FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3952" *)
  wire FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3968" *)
  wire FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3984" *)
  wire FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2360" *)
  wire [48:0] FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2351" *)
  wire [48:0] FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2354" *)
  wire [48:0] FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2357" *)
  wire [48:0] FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1395" *)
  reg [49:0] FpAdd_8U_23U_2_int_mant_p1_1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1363" *)
  reg [49:0] FpAdd_8U_23U_2_int_mant_p1_2_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1331" *)
  reg [49:0] FpAdd_8U_23U_2_int_mant_p1_3_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1299" *)
  reg [49:0] FpAdd_8U_23U_2_int_mant_p1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1902" *)
  wire FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1903" *)
  wire FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1904" *)
  wire FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2500" *)
  wire FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2617" *)
  wire FpAdd_8U_23U_2_is_a_greater_acc_1_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3913" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpAdd_8U_23U_2_is_a_greater_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2618" *)
  wire FpAdd_8U_23U_2_is_a_greater_acc_2_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3915" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpAdd_8U_23U_2_is_a_greater_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2619" *)
  wire FpAdd_8U_23U_2_is_a_greater_acc_3_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3917" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpAdd_8U_23U_2_is_a_greater_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2616" *)
  wire FpAdd_8U_23U_2_is_a_greater_acc_itm_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3911" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] FpAdd_8U_23U_2_is_a_greater_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1462" *)
  reg FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1492" *)
  reg FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1522" *)
  reg FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1552" *)
  reg FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2525" *)
  wire FpAdd_8U_23U_2_is_a_greater_oelse_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2665" *)
  wire FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4183" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2666" *)
  wire FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4185" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2667" *)
  wire FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4187" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2664" *)
  wire FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4181" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2473" *)
  wire FpAdd_8U_23U_2_is_addition_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1769" *)
  wire FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1466" *)
  reg FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1765" *)
  wire FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1496" *)
  reg FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1761" *)
  wire FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1526" *)
  reg FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2575" *)
  wire FpAdd_8U_23U_2_is_inf_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1757" *)
  wire FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1556" *)
  reg FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1589" *)
  reg FpAdd_8U_23U_2_mux_13_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1590" *)
  reg FpAdd_8U_23U_2_mux_13_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1614" *)
  reg FpAdd_8U_23U_2_mux_17_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1588" *)
  reg FpAdd_8U_23U_2_mux_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1615" *)
  reg FpAdd_8U_23U_2_mux_29_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1616" *)
  reg FpAdd_8U_23U_2_mux_29_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1642" *)
  reg FpAdd_8U_23U_2_mux_33_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1643" *)
  reg FpAdd_8U_23U_2_mux_45_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1644" *)
  reg FpAdd_8U_23U_2_mux_45_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1673" *)
  reg FpAdd_8U_23U_2_mux_49_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1674" *)
  reg FpAdd_8U_23U_2_mux_61_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1675" *)
  reg FpAdd_8U_23U_2_mux_61_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1465" *)
  reg [7:0] FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1495" *)
  reg [7:0] FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1525" *)
  reg [7:0] FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1991" *)
  wire FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1996" *)
  wire FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2002" *)
  wire FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1985" *)
  wire FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1555" *)
  reg [7:0] FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2233" *)
  wire [22:0] FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1471" *)
  reg [22:0] FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2235" *)
  wire [22:0] FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1501" *)
  reg [22:0] FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2237" *)
  wire [22:0] FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1531" *)
  reg [22:0] FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2239" *)
  wire [22:0] FpAdd_8U_23U_2_o_mant_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1561" *)
  reg [22:0] FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1463" *)
  reg [7:0] FpAdd_8U_23U_2_qr_2_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1464" *)
  reg [7:0] FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1493" *)
  reg [7:0] FpAdd_8U_23U_2_qr_3_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1494" *)
  reg [7:0] FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1523" *)
  reg [7:0] FpAdd_8U_23U_2_qr_4_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1524" *)
  reg [7:0] FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1553" *)
  reg [7:0] FpAdd_8U_23U_2_qr_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1554" *)
  reg [7:0] FpAdd_8U_23U_2_qr_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1049" *)
  wire [7:0] FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3887" *)
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3893" *)
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3899" *)
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3905" *)
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2288" *)
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2304" *)
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2320" *)
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2336" *)
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3291" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3292" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3275" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3276" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3283" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3284" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3267" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3268" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qelse_mux_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2290" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2306" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2322" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2338" *)
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2301" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_13_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2285" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_19_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2333" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_1_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2317" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_7_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2286" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2302" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2318" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2334" *)
  wire [48:0] FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2287" *)
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2303" *)
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2319" *)
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2335" *)
  wire [48:0] FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3933" *)
  wire FpAdd_8U_23U_and_35_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3949" *)
  wire FpAdd_8U_23U_and_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3965" *)
  wire FpAdd_8U_23U_and_39_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3981" *)
  wire FpAdd_8U_23U_and_41_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2432" *)
  wire FpAdd_8U_23U_and_43_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2425" *)
  wire FpAdd_8U_23U_and_45_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2418" *)
  wire FpAdd_8U_23U_and_47_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2411" *)
  wire FpAdd_8U_23U_and_49_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2431" *)
  wire FpAdd_8U_23U_and_51_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2424" *)
  wire FpAdd_8U_23U_and_53_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2417" *)
  wire FpAdd_8U_23U_and_55_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2410" *)
  wire FpAdd_8U_23U_and_57_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3930" *)
  wire FpAdd_8U_23U_and_59_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3931" *)
  wire FpAdd_8U_23U_and_61_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3946" *)
  wire FpAdd_8U_23U_and_63_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3947" *)
  wire FpAdd_8U_23U_and_65_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3962" *)
  wire FpAdd_8U_23U_and_67_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3963" *)
  wire FpAdd_8U_23U_and_69_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3978" *)
  wire FpAdd_8U_23U_and_71_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3979" *)
  wire FpAdd_8U_23U_and_73_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1945" *)
  wire [22:0] FpAdd_8U_23U_asn_35_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1944" *)
  wire [22:0] FpAdd_8U_23U_asn_40_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1943" *)
  wire [22:0] FpAdd_8U_23U_asn_45_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2223" *)
  wire [22:0] FpAdd_8U_23U_asn_50_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2169" *)
  wire FpAdd_8U_23U_b_right_shift_qif_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2172" *)
  wire FpAdd_8U_23U_b_right_shift_qif_and_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2173" *)
  wire FpAdd_8U_23U_b_right_shift_qif_and_tmp_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2176" *)
  wire FpAdd_8U_23U_b_right_shift_qif_and_tmp_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2289" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2305" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2321" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2337" *)
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3927" *)
  wire FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3943" *)
  wire FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3959" *)
  wire FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3975" *)
  wire FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2358" *)
  wire [48:0] FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2349" *)
  wire [48:0] FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2352" *)
  wire [48:0] FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2355" *)
  wire [48:0] FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2655" *)
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4097" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2652" *)
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4091" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2653" *)
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4093" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2654" *)
  wire FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_itm_23_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4095" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22" *)
  wire [23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1771" *)
  wire FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1767" *)
  wire FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1763" *)
  wire FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1759" *)
  wire FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1831" *)
  wire [7:0] FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1830" *)
  wire [7:0] FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2416" *)
  wire FpAdd_8U_23U_o_expo_and_1_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2423" *)
  wire FpAdd_8U_23U_o_expo_and_2_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2430" *)
  wire FpAdd_8U_23U_o_expo_and_3_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2409" *)
  wire FpAdd_8U_23U_o_expo_and_ssc;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1829" *)
  wire [7:0] FpAdd_8U_23U_o_expo_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2954" *)
  wire FpAdd_8U_23U_o_expo_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2905" *)
  wire FpAdd_8U_23U_o_expo_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2847" *)
  wire FpAdd_8U_23U_o_expo_or_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3004" *)
  wire FpAdd_8U_23U_o_expo_or_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2231" *)
  wire [22:0] FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1828" *)
  wire [22:0] FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1827" *)
  wire [22:0] FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1826" *)
  wire [22:0] FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1751" *)
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_2_itm_1_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1753" *)
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_3_itm_1_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1755" *)
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_4_itm_1_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1749" *)
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_itm_1_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3515" *)
  wire [7:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2462" *)
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2464" *)
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2466" *)
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2459" *)
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1472" *)
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1502" *)
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1532" *)
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1562" *)
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4020" *)
  wire [8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4031" *)
  wire [8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4042" *)
  wire [8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4009" *)
  wire [8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1750" *)
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_2_itm_1_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1752" *)
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_3_itm_1_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1754" *)
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_4_itm_1_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1748" *)
  reg FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_1_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1941" *)
  wire [7:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2461" *)
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2463" *)
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2465" *)
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2458" *)
  wire FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1455" *)
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1486" *)
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1516" *)
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1546" *)
  reg [255:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4015" *)
  wire [8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4026" *)
  wire [8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4037" *)
  wire [8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4004" *)
  wire [8:0] FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2559" *)
  wire FpMantRNE_49U_24U_1_else_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1453" *)
  reg FpMantRNE_49U_24U_1_else_carry_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2182" *)
  wire FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1484" *)
  reg FpMantRNE_49U_24U_1_else_carry_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2184" *)
  wire FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1514" *)
  reg FpMantRNE_49U_24U_1_else_carry_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2186" *)
  wire FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1544" *)
  reg FpMantRNE_49U_24U_1_else_carry_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2188" *)
  wire FpMantRNE_49U_24U_1_else_carry_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2447" *)
  wire FpMantRNE_49U_24U_1_else_o_mant_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2452" *)
  wire FpMantRNE_49U_24U_1_else_o_mant_and_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2455" *)
  wire FpMantRNE_49U_24U_1_else_o_mant_and_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2441" *)
  wire FpMantRNE_49U_24U_1_else_o_mant_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1467" *)
  reg FpMantRNE_49U_24U_2_else_carry_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2183" *)
  wire FpMantRNE_49U_24U_2_else_carry_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1497" *)
  reg FpMantRNE_49U_24U_2_else_carry_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2185" *)
  wire FpMantRNE_49U_24U_2_else_carry_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1527" *)
  reg FpMantRNE_49U_24U_2_else_carry_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2187" *)
  wire FpMantRNE_49U_24U_2_else_carry_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2446" *)
  wire FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1557" *)
  reg FpMantRNE_49U_24U_2_else_carry_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2189" *)
  wire FpMantRNE_49U_24U_2_else_carry_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4053" *)
  wire [48:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2925" *)
  wire [7:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4057" *)
  wire [48:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2975" *)
  wire [7:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4061" *)
  wire [48:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3025" *)
  wire [7:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4065" *)
  wire [48:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2869" *)
  wire [7:0] FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2368" *)
  wire FpNormalize_8U_49U_2_oelse_not_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2370" *)
  wire FpNormalize_8U_49U_2_oelse_not_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2372" *)
  wire FpNormalize_8U_49U_2_oelse_not_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2366" *)
  wire FpNormalize_8U_49U_2_oelse_not_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2904" *)
  wire [5:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2846" *)
  wire [5:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4051" *)
  wire [48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2903" *)
  wire [1:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4055" *)
  wire [48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2951" *)
  wire [1:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4059" *)
  wire [48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3001" *)
  wire [1:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4063" *)
  wire [48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3003" *)
  wire [5:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2953" *)
  wire [5:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2845" *)
  wire [1:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2367" *)
  wire FpNormalize_8U_49U_oelse_not_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2369" *)
  wire FpNormalize_8U_49U_oelse_not_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2371" *)
  wire FpNormalize_8U_49U_oelse_not_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2365" *)
  wire FpNormalize_8U_49U_oelse_not_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1911" *)
  wire [30:0] IntLog2_32U_IntLog2_32U_mux_1_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1913" *)
  wire [30:0] IntLog2_32U_IntLog2_32U_mux_2_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1909" *)
  wire [30:0] IntLog2_32U_IntLog2_32U_mux_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1233" *)
  reg [30:0] IntLog2_32U_ac_int_cctor_1_30_0_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1234" *)
  reg [30:0] IntLog2_32U_ac_int_cctor_1_30_0_2_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1235" *)
  reg [30:0] IntLog2_32U_ac_int_cctor_1_30_0_3_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1236" *)
  reg [30:0] IntLog2_32U_ac_int_cctor_1_30_0_sva_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2112" *)
  wire [30:0] IntLog2_32U_mux1h_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2350" *)
  wire [8:0] IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2353" *)
  wire [8:0] IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2356" *)
  wire [8:0] IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2359" *)
  wire [8:0] IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1473" *)
  reg IsNaN_8U_23U_10_land_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1474" *)
  reg IsNaN_8U_23U_10_land_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1503" *)
  reg IsNaN_8U_23U_10_land_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1504" *)
  reg IsNaN_8U_23U_10_land_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1533" *)
  reg IsNaN_8U_23U_10_land_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1534" *)
  reg IsNaN_8U_23U_10_land_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1563" *)
  reg IsNaN_8U_23U_10_land_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1564" *)
  reg IsNaN_8U_23U_10_land_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2544" *)
  wire IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2491" *)
  wire IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_3_aelse_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2537" *)
  wire IsNaN_8U_23U_1_aelse_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2536" *)
  wire IsNaN_8U_23U_1_aelse_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1266" *)
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1267" *)
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1268" *)
  reg IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1259" *)
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1260" *)
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1261" *)
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2230" *)
  wire IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1253" *)
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1254" *)
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1246" *)
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1247" *)
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1248" *)
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2533" *)
  wire IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2483" *)
  wire IsNaN_8U_23U_3_aelse_and_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2443" *)
  wire IsNaN_8U_23U_3_aelse_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1454" *)
  reg IsNaN_8U_23U_3_land_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2179" *)
  wire IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1693" *)
  reg IsNaN_8U_23U_3_land_1_lpi_1_dfm_st_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1485" *)
  reg IsNaN_8U_23U_3_land_2_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1705" *)
  reg IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1706" *)
  reg IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1515" *)
  reg IsNaN_8U_23U_3_land_3_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1716" *)
  reg IsNaN_8U_23U_3_land_3_lpi_1_dfm_st_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1545" *)
  reg IsNaN_8U_23U_3_land_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1907" *)
  wire IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1729" *)
  reg IsNaN_8U_23U_3_land_lpi_1_dfm_st_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1031" *)
  wire IsNaN_8U_23U_3_nor_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1034" *)
  wire IsNaN_8U_23U_3_nor_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1028" *)
  wire IsNaN_8U_23U_3_nor_6_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1037" *)
  wire IsNaN_8U_23U_3_nor_8_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1658" *)
  reg IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1576" *)
  reg IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1806" *)
  wire IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1265" *)
  reg IsNaN_8U_23U_4_land_1_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2209" *)
  wire IsNaN_8U_23U_4_land_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1258" *)
  reg IsNaN_8U_23U_4_land_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1252" *)
  reg IsNaN_8U_23U_4_land_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1245" *)
  reg IsNaN_8U_23U_4_land_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2208" *)
  wire IsNaN_8U_23U_4_land_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1657" *)
  reg IsNaN_8U_23U_4_nor_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1575" *)
  reg IsNaN_8U_23U_4_nor_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1080" *)
  wire IsNaN_8U_23U_4_nor_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1047" *)
  wire IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1044" *)
  wire IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1041" *)
  wire IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2566" *)
  wire IsNaN_8U_23U_5_IsNaN_8U_23U_6_aelse_or_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1456" *)
  reg IsNaN_8U_23U_6_land_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1457" *)
  reg IsNaN_8U_23U_6_land_1_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1487" *)
  reg IsNaN_8U_23U_6_land_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1488" *)
  reg IsNaN_8U_23U_6_land_2_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1517" *)
  reg IsNaN_8U_23U_6_land_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1518" *)
  reg IsNaN_8U_23U_6_land_3_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1547" *)
  reg IsNaN_8U_23U_6_land_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1548" *)
  reg IsNaN_8U_23U_6_land_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2548" *)
  wire IsNaN_8U_23U_7_aelse_and_17_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1469" *)
  reg IsNaN_8U_23U_7_land_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1470" *)
  reg IsNaN_8U_23U_7_land_1_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1697" *)
  reg IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1698" *)
  reg IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1699" *)
  reg IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1499" *)
  reg IsNaN_8U_23U_7_land_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1500" *)
  reg IsNaN_8U_23U_7_land_2_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1709" *)
  reg IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1710" *)
  reg IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1529" *)
  reg IsNaN_8U_23U_7_land_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1530" *)
  reg IsNaN_8U_23U_7_land_3_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1719" *)
  reg IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1720" *)
  reg IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1721" *)
  reg IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1559" *)
  reg IsNaN_8U_23U_7_land_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1560" *)
  reg IsNaN_8U_23U_7_land_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1732" *)
  reg IsNaN_8U_23U_7_land_lpi_1_dfm_st_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1640" *)
  reg IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1805" *)
  wire IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1671" *)
  reg IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2451" *)
  wire IsNaN_8U_23U_8_aelse_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2490" *)
  wire IsNaN_8U_23U_8_and_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2489" *)
  wire IsNaN_8U_23U_8_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1262" *)
  reg IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1255" *)
  reg IsNaN_8U_23U_8_land_2_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1256" *)
  reg IsNaN_8U_23U_8_land_2_lpi_1_dfm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1249" *)
  reg IsNaN_8U_23U_8_land_3_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1250" *)
  reg IsNaN_8U_23U_8_land_3_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1242" *)
  reg IsNaN_8U_23U_8_land_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1243" *)
  reg IsNaN_8U_23U_8_land_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1639" *)
  reg IsNaN_8U_23U_8_nor_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1079" *)
  wire IsNaN_8U_23U_8_nor_2_tmp_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1670" *)
  reg IsNaN_8U_23U_8_nor_3_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2478" *)
  wire IsZero_8U_23U_1_IsZero_8U_23U_4_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2517" *)
  wire IsZero_8U_23U_4_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2476" *)
  wire IsZero_8U_23U_4_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1040" *)
  wire IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1050" *)
  wire IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1046" *)
  wire IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1043" *)
  wire IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2481" *)
  wire IsZero_8U_23U_7_and_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1045" *)
  wire IsZero_8U_23U_8_IsZero_8U_23U_8_nor_1_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1042" *)
  wire IsZero_8U_23U_8_IsZero_8U_23U_8_nor_2_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1039" *)
  wire IsZero_8U_23U_8_IsZero_8U_23U_8_nor_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1048" *)
  wire IsZero_8U_23U_8_IsZero_8U_23U_8_nor_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3277" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3281" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3265" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3293" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3269" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3289" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3273" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3285" *)
  (* unused_bits = "0" *)
  wire [8:0] acc_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3345" *)
  wire and_100_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3346" *)
  wire and_101_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3348" *)
  wire and_102_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3349" *)
  wire and_103_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3351" *)
  wire and_104_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3352" *)
  wire and_105_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3354" *)
  wire and_106_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3571" *)
  wire and_1089_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3356" *)
  wire and_108_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3357" *)
  wire and_109_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3359" *)
  wire and_110_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3360" *)
  wire and_111_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3362" *)
  wire and_112_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2494" *)
  wire and_1138_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2495" *)
  wire and_1139_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3368" *)
  wire and_113_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2496" *)
  wire and_1140_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2497" *)
  wire and_1141_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2492" *)
  wire and_1142_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3724" *)
  wire and_1146_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3692" *)
  wire and_1147_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3714" *)
  wire and_1148_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3704" *)
  wire and_1149_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3380" *)
  wire and_114_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3640" *)
  wire and_1151_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3632" *)
  wire and_1153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3583" *)
  wire and_1156_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3576" *)
  wire and_1158_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3386" *)
  wire and_115_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3532" *)
  wire and_1160_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3525" *)
  wire and_1162_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3459" *)
  wire and_1164_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3451" *)
  wire and_1166_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3394" *)
  wire and_116_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3647" *)
  wire and_1174_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3628" *)
  wire and_1176_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3702" *)
  wire and_1179_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3400" *)
  wire and_117_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3408" *)
  wire and_118_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3414" *)
  wire and_119_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3424" *)
  wire and_120_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3461" *)
  wire and_127_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3489" *)
  wire and_131_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3503" *)
  wire and_132_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2573" *)
  wire and_134_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3534" *)
  wire and_138_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3547" *)
  wire and_142_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3559" *)
  wire and_143_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3573" *)
  wire and_147_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3585" *)
  wire and_149_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3598" *)
  wire and_152_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3610" *)
  wire and_153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3623" *)
  wire and_158_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3642" *)
  wire and_160_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3659" *)
  wire and_163_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3671" *)
  wire and_164_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3674" *)
  wire and_166_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2580" *)
  wire and_178_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3694" *)
  wire and_179_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3706" *)
  wire and_193_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3716" *)
  wire and_204_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3726" *)
  wire and_215_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3780" *)
  wire and_219_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3783" *)
  wire and_220_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3786" *)
  wire and_221_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3792" *)
  wire and_222_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3795" *)
  wire and_224_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3797" *)
  wire and_226_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3803" *)
  wire and_228_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3806" *)
  wire and_230_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3808" *)
  wire and_232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3814" *)
  wire and_233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3817" *)
  wire and_235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3820" *)
  wire and_236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1960" *)
  wire and_284_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1961" *)
  wire and_286_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1962" *)
  wire and_288_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1963" *)
  wire and_290_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1964" *)
  wire and_292_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1965" *)
  wire and_300_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1966" *)
  wire and_302_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1967" *)
  wire and_304_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1968" *)
  wire and_306_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1969" *)
  wire and_308_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1970" *)
  wire and_316_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1971" *)
  wire and_318_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1972" *)
  wire and_320_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1973" *)
  wire and_322_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1974" *)
  wire and_324_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1975" *)
  wire and_330_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1976" *)
  wire and_332_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1977" *)
  wire and_334_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1978" *)
  wire and_336_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1979" *)
  wire and_338_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1980" *)
  wire and_344_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1981" *)
  wire and_347_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1843" *)
  wire and_355_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1988" *)
  wire and_364_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1842" *)
  wire and_375_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2534" *)
  wire and_401_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2546" *)
  wire and_427_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2005" *)
  wire and_428_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2540" *)
  wire and_42_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2006" *)
  wire and_430_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3127" *)
  wire and_447_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3157" *)
  wire and_451_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3189" *)
  wire and_455_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3218" *)
  wire and_459_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2865" *)
  wire and_45_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1862" *)
  wire and_465_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1863" *)
  wire and_466_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2921" *)
  wire and_48_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2932" *)
  wire and_49_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2007" *)
  wire and_524_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2008" *)
  wire and_525_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2009" *)
  wire and_527_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2010" *)
  wire and_529_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2971" *)
  wire and_54_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2011" *)
  wire and_551_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1840" *)
  wire and_553_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1841" *)
  wire and_555_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2014" *)
  wire and_559_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1839" *)
  wire and_562_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2017" *)
  wire and_564_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2018" *)
  wire and_566_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1838" *)
  wire and_567_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2021" *)
  wire and_570_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1837" *)
  wire and_572_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2024" *)
  wire and_574_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2025" *)
  wire and_576_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1836" *)
  wire and_577_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2028" *)
  wire and_580_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1835" *)
  wire and_582_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2031" *)
  wire and_586_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2032" *)
  wire and_588_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1833" *)
  wire and_590_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1834" *)
  wire and_592_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2035" *)
  wire and_595_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1832" *)
  wire and_597_m1c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3021" *)
  wire and_59_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2038" *)
  wire and_604_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2039" *)
  wire and_606_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3056" *)
  wire and_62_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2550" *)
  wire and_636_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3061" *)
  wire and_63_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3477" *)
  wire and_649_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3062" *)
  wire and_64_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2041" *)
  wire and_653_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3542" *)
  wire and_657_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2044" *)
  wire and_661_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3593" *)
  wire and_665_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2047" *)
  wire and_668_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3654" *)
  wire and_672_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2049" *)
  wire and_676_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2051" *)
  wire and_679_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3078" *)
  wire and_69_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3082" *)
  wire and_70_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3083" *)
  wire and_71_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3099" *)
  wire and_74_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3102" *)
  wire and_75_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3103" *)
  wire and_76_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3836" *)
  wire and_773_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3832" *)
  wire and_774_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1879" *)
  wire and_780_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1877" *)
  wire and_784_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1876" *)
  wire and_787_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1875" *)
  wire and_789_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1878" *)
  wire and_794_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1874" *)
  wire and_795_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3119" *)
  wire and_79_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3645" *)
  wire and_804_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3588" *)
  wire and_808_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3123" *)
  wire and_80_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1872" *)
  wire and_811_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3537" *)
  wire and_812_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1871" *)
  wire and_814_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3486" *)
  wire and_815_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3487" *)
  wire and_816_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3464" *)
  wire and_819_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3124" *)
  wire and_81_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3432" *)
  wire and_822_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3426" *)
  wire and_823_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2557" *)
  wire and_826_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3340" *)
  wire and_827_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1855" *)
  wire and_82_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3263" *)
  wire and_830_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2541" *)
  wire and_832_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1857" *)
  wire and_835_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1856" *)
  wire and_839_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2583" *)
  wire and_843_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1854" *)
  wire and_846_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1893" *)
  wire and_848_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1892" *)
  wire and_850_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2564" *)
  wire and_852_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1853" *)
  wire and_854_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3011" *)
  wire and_858_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3013" *)
  wire and_859_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2961" *)
  wire and_861_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2963" *)
  wire and_862_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2911" *)
  wire and_864_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2913" *)
  wire and_865_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2855" *)
  wire and_868_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2857" *)
  wire and_869_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1947" *)
  wire and_896_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2553" *)
  wire and_898_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2554" *)
  wire and_901_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1950" *)
  wire and_905_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2555" *)
  wire and_907_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2506" *)
  wire and_956_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2507" *)
  wire and_961_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3342" *)
  wire and_98_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1197" *)
  wire and_dcpl_148;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1199" *)
  wire and_dcpl_161;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1200" *)
  wire and_dcpl_162;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1214" *)
  wire and_dcpl_258;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1215" *)
  wire and_dcpl_259;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1216" *)
  wire and_dcpl_280;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1217" *)
  wire and_dcpl_284;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1218" *)
  wire and_dcpl_288;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1219" *)
  wire and_dcpl_292;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1220" *)
  wire and_dcpl_296;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1221" *)
  wire and_dcpl_300;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1222" *)
  wire and_dcpl_304;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1223" *)
  wire and_dcpl_308;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1224" *)
  wire and_dcpl_309;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1225" *)
  wire and_dcpl_314;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1226" *)
  wire and_dcpl_315;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1227" *)
  wire and_dcpl_316;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1228" *)
  wire and_dcpl_351;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1229" *)
  wire and_dcpl_364;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1230" *)
  wire and_dcpl_403;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1231" *)
  wire and_dcpl_405;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1188" *)
  wire and_dcpl_54;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1959" *)
  wire and_dcpl_540;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1983" *)
  wire and_dcpl_576;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1189" *)
  wire and_dcpl_59;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1190" *)
  wire and_dcpl_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2040" *)
  wire and_dcpl_648;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1191" *)
  wire and_dcpl_67;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1192" *)
  wire and_dcpl_71;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1193" *)
  wire and_dcpl_72;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1194" *)
  wire and_dcpl_74;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1196" *)
  wire and_dcpl_98;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3323" *)
  wire and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1169" *)
  wire and_tmp_103;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1172" *)
  wire and_tmp_108;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1173" *)
  wire and_tmp_113;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1176" *)
  wire and_tmp_119;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1177" *)
  wire and_tmp_124;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1178" *)
  wire and_tmp_130;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1180" *)
  wire and_tmp_131;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1104" *)
  wire and_tmp_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1187" *)
  wire and_tmp_178;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1107" *)
  wire and_tmp_19;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2159" *)
  wire and_tmp_201;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1115" *)
  wire and_tmp_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1089" *)
  wire and_tmp_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1155" *)
  wire and_tmp_59;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1090" *)
  wire and_tmp_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1156" *)
  wire and_tmp_61;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1158" *)
  wire and_tmp_69;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1160" *)
  wire and_tmp_83;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1164" *)
  wire and_tmp_92;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1166" *)
  wire and_tmp_97;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1168" *)
  wire and_tmp_98;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1443" *)
  reg cfg_lut_hybrid_priority_1_sva_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1439" *)
  reg cfg_lut_hybrid_priority_1_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1440" *)
  reg cfg_lut_hybrid_priority_1_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1441" *)
  reg cfg_lut_hybrid_priority_1_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1442" *)
  reg cfg_lut_hybrid_priority_1_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2467" *)
  wire cfg_lut_hybrid_priority_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:951" *)
  input cfg_lut_hybrid_priority_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:976" *)
  wire cfg_lut_hybrid_priority_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1428" *)
  reg cfg_lut_le_function_1_sva_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1724" *)
  reg cfg_lut_le_function_1_sva_st_41;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1725" *)
  reg cfg_lut_le_function_1_sva_st_42;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:948" *)
  input cfg_lut_le_function_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:973" *)
  wire cfg_lut_le_function_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1418" *)
  reg [7:0] cfg_lut_le_index_offset_1_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1419" *)
  reg [7:0] cfg_lut_le_index_offset_1_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1420" *)
  reg [7:0] cfg_lut_le_index_offset_1_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1421" *)
  reg [7:0] cfg_lut_le_index_offset_1_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2434" *)
  wire cfg_lut_le_index_offset_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:945" *)
  input [7:0] cfg_lut_le_index_offset_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:970" *)
  wire [7:0] cfg_lut_le_index_offset_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1422" *)
  reg [7:0] cfg_lut_le_index_select_1_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1423" *)
  reg [7:0] cfg_lut_le_index_select_1_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1424" *)
  reg [7:0] cfg_lut_le_index_select_1_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:946" *)
  input [7:0] cfg_lut_le_index_select_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:971" *)
  wire [7:0] cfg_lut_le_index_select_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1740" *)
  reg [30:0] cfg_lut_le_start_1_sva_2_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1741" *)
  reg [30:0] cfg_lut_le_start_1_sva_3_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1416" *)
  reg [31:0] cfg_lut_le_start_1_sva_41;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2440" *)
  wire cfg_lut_le_start_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:943" *)
  input [31:0] cfg_lut_le_start_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:968" *)
  wire [31:0] cfg_lut_le_start_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1425" *)
  reg [7:0] cfg_lut_lo_index_select_1_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1426" *)
  reg [7:0] cfg_lut_lo_index_select_1_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1427" *)
  reg [7:0] cfg_lut_lo_index_select_1_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:947" *)
  input [7:0] cfg_lut_lo_index_select_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:972" *)
  wire [7:0] cfg_lut_lo_index_select_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1742" *)
  reg [30:0] cfg_lut_lo_start_1_sva_2_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1743" *)
  reg [30:0] cfg_lut_lo_start_1_sva_3_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1417" *)
  reg [31:0] cfg_lut_lo_start_1_sva_41;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:944" *)
  input [31:0] cfg_lut_lo_start_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:969" *)
  wire [31:0] cfg_lut_lo_start_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1438" *)
  reg cfg_lut_oflow_priority_1_sva_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1434" *)
  reg cfg_lut_oflow_priority_1_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1435" *)
  reg cfg_lut_oflow_priority_1_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1436" *)
  reg cfg_lut_oflow_priority_1_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1437" *)
  reg cfg_lut_oflow_priority_1_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:950" *)
  input cfg_lut_oflow_priority_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:975" *)
  wire cfg_lut_oflow_priority_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1433" *)
  reg cfg_lut_uflow_priority_1_sva_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1429" *)
  reg cfg_lut_uflow_priority_1_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1430" *)
  reg cfg_lut_uflow_priority_1_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1431" *)
  reg cfg_lut_uflow_priority_1_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1432" *)
  reg cfg_lut_uflow_priority_1_sva_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:949" *)
  input cfg_lut_uflow_priority_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:974" *)
  wire cfg_lut_uflow_priority_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1444" *)
  reg [1:0] cfg_precision_1_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1733" *)
  reg [1:0] cfg_precision_1_sva_st_107;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1688" *)
  reg [1:0] cfg_precision_1_sva_st_70;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1689" *)
  reg [1:0] cfg_precision_1_sva_st_71;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1694" *)
  reg [1:0] cfg_precision_1_sva_st_72;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2460" *)
  wire cfg_precision_and_24_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2433" *)
  wire cfg_precision_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:952" *)
  input [1:0] cfg_precision_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:977" *)
  wire [1:0] cfg_precision_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:942" *)
  output chn_lut_in_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:941" *)
  input chn_lut_in_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:940" *)
  input [127:0] chn_lut_in_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:963" *)
  wire chn_lut_in_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:966" *)
  wire [127:0] chn_lut_in_rsci_d_mxwt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:962" *)
  reg chn_lut_in_rsci_iswt0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:965" *)
  reg chn_lut_in_rsci_ld_core_psct;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2177" *)
  wire chn_lut_in_rsci_ld_core_psct_mx0c0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:956" *)
  input chn_lut_in_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:957" *)
  output chn_lut_in_rsci_oswt_unreg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:964" *)
  wire chn_lut_in_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1845" *)
  wire chn_lut_out_and_13_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1846" *)
  wire chn_lut_out_and_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1847" *)
  wire chn_lut_out_and_15_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1848" *)
  wire chn_lut_out_and_16_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1844" *)
  wire chn_lut_out_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:955" *)
  output chn_lut_out_rsc_lz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:954" *)
  input chn_lut_out_rsc_vz;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:953" *)
  output [323:0] chn_lut_out_rsc_z;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:979" *)
  wire chn_lut_out_rsci_bawt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1020" *)
  reg [22:0] chn_lut_out_rsci_d_104_82;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1019" *)
  reg [11:0] chn_lut_out_rsci_d_116_105;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1025" *)
  reg [11:0] chn_lut_out_rsci_d_11_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1018" *)
  reg [22:0] chn_lut_out_rsci_d_139_117;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1017" *)
  reg [127:0] chn_lut_out_rsci_d_267_140;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1016" *)
  reg chn_lut_out_rsci_d_268;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1015" *)
  reg chn_lut_out_rsci_d_269;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1014" *)
  reg chn_lut_out_rsci_d_270;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1013" *)
  reg chn_lut_out_rsci_d_271;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1012" *)
  reg chn_lut_out_rsci_d_272;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1011" *)
  reg chn_lut_out_rsci_d_273;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1010" *)
  reg chn_lut_out_rsci_d_274;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1009" *)
  reg chn_lut_out_rsci_d_275;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1008" *)
  reg chn_lut_out_rsci_d_276;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1007" *)
  reg chn_lut_out_rsci_d_277;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1006" *)
  reg chn_lut_out_rsci_d_278;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1005" *)
  reg chn_lut_out_rsci_d_279;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1004" *)
  reg [5:0] chn_lut_out_rsci_d_285_280;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1003" *)
  reg chn_lut_out_rsci_d_286;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1002" *)
  reg chn_lut_out_rsci_d_287;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1001" *)
  reg chn_lut_out_rsci_d_288;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1000" *)
  reg [5:0] chn_lut_out_rsci_d_294_289;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:999" *)
  reg chn_lut_out_rsci_d_295;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:998" *)
  reg chn_lut_out_rsci_d_296;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:997" *)
  reg chn_lut_out_rsci_d_297;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:996" *)
  reg [5:0] chn_lut_out_rsci_d_303_298;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:995" *)
  reg chn_lut_out_rsci_d_304;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:994" *)
  reg chn_lut_out_rsci_d_305;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:993" *)
  reg chn_lut_out_rsci_d_306;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:992" *)
  reg [5:0] chn_lut_out_rsci_d_312_307;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:991" *)
  reg chn_lut_out_rsci_d_313;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:990" *)
  reg chn_lut_out_rsci_d_314;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:989" *)
  reg chn_lut_out_rsci_d_315;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:988" *)
  reg chn_lut_out_rsci_d_316;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:987" *)
  reg chn_lut_out_rsci_d_317;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:986" *)
  reg chn_lut_out_rsci_d_318;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:985" *)
  reg chn_lut_out_rsci_d_319;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:984" *)
  reg chn_lut_out_rsci_d_320;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:983" *)
  reg chn_lut_out_rsci_d_321;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:982" *)
  reg chn_lut_out_rsci_d_322;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:981" *)
  reg chn_lut_out_rsci_d_323;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1024" *)
  reg [22:0] chn_lut_out_rsci_d_34_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1023" *)
  reg [11:0] chn_lut_out_rsci_d_46_35;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1022" *)
  reg [22:0] chn_lut_out_rsci_d_69_47;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1021" *)
  reg [11:0] chn_lut_out_rsci_d_81_70;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:978" *)
  reg chn_lut_out_rsci_iswt0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:958" *)
  input chn_lut_out_rsci_oswt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:959" *)
  output chn_lut_out_rsci_oswt_unreg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:980" *)
  wire chn_lut_out_rsci_wen_comp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:961" *)
  wire core_wen;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:967" *)
  wire core_wten;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1026" *)
  wire [1:0] fsm_output;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2393" *)
  wire [5:0] libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2394" *)
  wire [5:0] libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2395" *)
  wire [5:0] libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2396" *)
  wire [5:0] libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2397" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2398" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2399" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2400" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2401" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2402" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_17;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2403" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_18;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2404" *)
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_19;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1445" *)
  reg [127:0] lut_in_data_sva_154;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1446" *)
  reg [127:0] lut_in_data_sva_155;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1447" *)
  reg [127:0] lut_in_data_sva_156;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1448" *)
  reg [127:0] lut_in_data_sva_157;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1449" *)
  reg [127:0] lut_in_data_sva_158;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1573" *)
  reg lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1574" *)
  reg lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2783" *)
  wire [49:0] lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2785" *)
  wire [49:0] lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2656" *)
  wire lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4115" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2660" *)
  wire lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4123" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1038" *)
  wire lut_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1586" *)
  reg lut_lookup_1_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4455" *)
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  wire [3:0] lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2793" *)
  wire [49:0] lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2791" *)
  wire [49:0] lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2620" *)
  wire lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3919" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2872" *)
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2624" *)
  wire lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3934" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3937" *)
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1036" *)
  wire lut_lookup_1_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2203" *)
  wire lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2204" *)
  wire lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2379" *)
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2377" *)
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2787" *)
  wire [49:0] lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2789" *)
  wire [49:0] lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2428" *)
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3928" *)
  wire [7:0] lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1591" *)
  reg [7:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2082" *)
  wire [34:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2633" *)
  wire lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4007" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246" *)
  wire [247:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1593" *)
  reg lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1063" *)
  wire [9:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2083" *)
  wire [255:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1581" *)
  reg [7:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2080" *)
  wire [34:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4005" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246" *)
  wire [247:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1582" *)
  reg lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1065" *)
  wire [9:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2081" *)
  wire [255:0] lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1577" *)
  reg [22:0] lut_lookup_1_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3891" *)
  wire [22:0] lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1468" *)
  reg lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1076" *)
  wire lut_lookup_1_FpMantRNE_49U_24U_2_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1587" *)
  reg [22:0] lut_lookup_1_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3888" *)
  wire [22:0] lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1078" *)
  wire lut_lookup_1_FpMantRNE_49U_24U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4099" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4101" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] lut_lookup_1_FpNormalize_8U_49U_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2870" *)
  wire [7:0] lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2130" *)
  wire [48:0] lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2426" *)
  wire [7:0] lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2128" *)
  wire [48:0] lut_lookup_1_FpNormalize_8U_49U_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3474" *)
  wire [30:0] lut_lookup_1_IntLog2_32U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3473" *)
  wire [30:0] lut_lookup_1_IntLog2_32U_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1571" *)
  reg [1:0] lut_lookup_1_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2113" *)
  wire [30:0] lut_lookup_1_IntLog2_32U_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2131" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126" *)
  wire [286:0] lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4054" *)
  wire lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1077" *)
  wire [8:0] lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2129" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126" *)
  wire [286:0] lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4052" *)
  wire lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1480" *)
  reg lut_lookup_1_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2612" *)
  wire lut_lookup_1_else_1_acc_itm_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3879" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_1_else_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3513" *)
  wire [8:0] lut_lookup_1_else_1_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2363" *)
  wire [31:0] lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1594" *)
  reg [31:0] lut_lookup_1_else_1_else_else_lo_data_f_and_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2145" *)
  wire [31:0] lut_lookup_1_else_1_else_else_lo_data_f_lshift_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2099" *)
  wire [34:0] lut_lookup_1_else_1_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1596" *)
  reg lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1597" *)
  reg lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1701" *)
  reg lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1595" *)
  reg lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1779" *)
  wire lut_lookup_1_else_2_and_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1778" *)
  wire lut_lookup_1_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2644" *)
  wire lut_lookup_1_else_else_acc_1_itm_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4075" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_1_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2224" *)
  wire [8:0] lut_lookup_1_else_else_else_else_acc_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2361" *)
  wire [31:0] lut_lookup_1_else_else_else_else_le_data_f_acc_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1583" *)
  reg [31:0] lut_lookup_1_else_else_else_else_le_data_f_and_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2144" *)
  wire [31:0] lut_lookup_1_else_else_else_else_le_data_f_lshift_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2098" *)
  wire [34:0] lut_lookup_1_else_else_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2597" *)
  wire lut_lookup_1_else_else_else_if_acc_itm_3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3845" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_1_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2632" *)
  wire lut_lookup_1_else_if_else_if_acc_itm_3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3999" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_1_else_if_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2596" *)
  wire lut_lookup_1_if_else_else_acc_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3843" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] lut_lookup_1_if_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2604" *)
  wire lut_lookup_1_if_else_else_else_else_acc_itm_32_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3859" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_1_if_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3492" *)
  wire [6:0] lut_lookup_1_if_else_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2097" *)
  wire [34:0] lut_lookup_1_if_else_else_else_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3494" *)
  wire [3:0] lut_lookup_1_if_else_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2096" *)
  wire [34:0] lut_lookup_1_if_else_else_else_else_if_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1692" *)
  reg lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1572" *)
  reg [5:0] lut_lookup_1_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2605" *)
  wire lut_lookup_1_if_else_else_else_if_acc_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3861" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_1_if_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1281" *)
  reg lut_lookup_1_if_else_slc_32_svs_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1282" *)
  reg lut_lookup_1_if_else_slc_32_svs_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1283" *)
  reg lut_lookup_1_if_else_slc_32_svs_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1284" *)
  reg lut_lookup_1_if_else_slc_32_svs_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1690" *)
  reg lut_lookup_1_if_else_slc_32_svs_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2628" *)
  wire lut_lookup_1_if_if_else_acc_itm_9_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3991" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8" *)
  wire [9:0] lut_lookup_1_if_if_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2640" *)
  wire lut_lookup_1_if_if_else_else_if_acc_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4067" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_1_if_if_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1601" *)
  reg lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1602" *)
  reg lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2795" *)
  wire [49:0] lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2797" *)
  wire [49:0] lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2657" *)
  wire lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4117" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2661" *)
  wire lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4125" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1035" *)
  wire lut_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1612" *)
  reg lut_lookup_2_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4501" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4490" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2805" *)
  wire [49:0] lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2803" *)
  wire [49:0] lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2621" *)
  wire lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3921" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2928" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2625" *)
  wire lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3950" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3953" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1033" *)
  wire lut_lookup_2_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2205" *)
  wire lut_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2383" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2381" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2799" *)
  wire [49:0] lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2801" *)
  wire [49:0] lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2421" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3944" *)
  wire [7:0] lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1617" *)
  reg [7:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2086" *)
  wire [34:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2635" *)
  wire lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4018" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246" *)
  wire [247:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1619" *)
  reg lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1059" *)
  wire [9:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2087" *)
  wire [255:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1607" *)
  reg [7:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2084" *)
  wire [34:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4016" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246" *)
  wire [247:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1608" *)
  reg lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1061" *)
  wire [9:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2085" *)
  wire [255:0] lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1603" *)
  reg [22:0] lut_lookup_2_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3897" *)
  wire [22:0] lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1498" *)
  reg lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1073" *)
  wire lut_lookup_2_FpMantRNE_49U_24U_2_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1613" *)
  reg [22:0] lut_lookup_2_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3894" *)
  wire [22:0] lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1075" *)
  wire lut_lookup_2_FpMantRNE_49U_24U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4103" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4105" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] lut_lookup_2_FpNormalize_8U_49U_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2926" *)
  wire [7:0] lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2134" *)
  wire [48:0] lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2419" *)
  wire [7:0] lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2132" *)
  wire [48:0] lut_lookup_2_FpNormalize_8U_49U_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3539" *)
  wire [30:0] lut_lookup_2_IntLog2_32U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3538" *)
  wire [30:0] lut_lookup_2_IntLog2_32U_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1599" *)
  reg [1:0] lut_lookup_2_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2119" *)
  wire [30:0] lut_lookup_2_IntLog2_32U_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2135" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126" *)
  wire [286:0] lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4058" *)
  wire lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1074" *)
  wire [8:0] lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2133" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126" *)
  wire [286:0] lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4056" *)
  wire lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1510" *)
  reg lut_lookup_2_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2613" *)
  wire lut_lookup_2_else_1_acc_itm_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3881" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_2_else_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1620" *)
  reg [31:0] lut_lookup_2_else_1_else_else_lo_data_f_and_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2103" *)
  wire [34:0] lut_lookup_2_else_1_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1622" *)
  reg lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1623" *)
  reg lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1712" *)
  reg lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1621" *)
  reg lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1782" *)
  wire lut_lookup_2_else_2_and_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1781" *)
  wire lut_lookup_2_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2646" *)
  wire lut_lookup_2_else_else_acc_1_itm_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4079" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_2_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1609" *)
  reg [31:0] lut_lookup_2_else_else_else_else_le_data_f_and_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2102" *)
  wire [34:0] lut_lookup_2_else_else_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2599" *)
  wire lut_lookup_2_else_else_else_if_acc_itm_3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3849" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_2_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2634" *)
  wire lut_lookup_2_else_if_else_if_acc_itm_3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4010" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_2_else_if_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2598" *)
  wire lut_lookup_2_if_else_else_acc_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3847" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] lut_lookup_2_if_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2606" *)
  wire lut_lookup_2_if_else_else_else_else_acc_itm_32_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3863" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_2_if_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3548" *)
  wire [6:0] lut_lookup_2_if_else_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2101" *)
  wire [34:0] lut_lookup_2_if_else_else_else_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3550" *)
  wire [3:0] lut_lookup_2_if_else_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2100" *)
  wire [34:0] lut_lookup_2_if_else_else_else_else_if_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1704" *)
  reg lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1600" *)
  reg [5:0] lut_lookup_2_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2607" *)
  wire lut_lookup_2_if_else_else_else_if_acc_itm_3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3865" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_2_if_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1277" *)
  reg lut_lookup_2_if_else_slc_32_svs_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1278" *)
  reg lut_lookup_2_if_else_slc_32_svs_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1279" *)
  reg lut_lookup_2_if_else_slc_32_svs_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1280" *)
  reg lut_lookup_2_if_else_slc_32_svs_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1702" *)
  reg lut_lookup_2_if_else_slc_32_svs_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2629" *)
  wire lut_lookup_2_if_if_else_acc_itm_9_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3993" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8" *)
  wire [9:0] lut_lookup_2_if_if_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2641" *)
  wire lut_lookup_2_if_if_else_else_if_acc_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4069" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_2_if_if_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1627" *)
  reg lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1628" *)
  reg lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2807" *)
  wire [49:0] lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2809" *)
  wire [49:0] lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2658" *)
  wire lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4119" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2662" *)
  wire lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4127" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1032" *)
  wire lut_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1638" *)
  reg lut_lookup_3_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4547" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4536" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2817" *)
  wire [49:0] lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2815" *)
  wire [49:0] lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2622" *)
  wire lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3923" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2978" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2626" *)
  wire lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3966" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3969" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1030" *)
  wire lut_lookup_3_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2206" *)
  wire lut_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2387" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2385" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2811" *)
  wire [49:0] lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2813" *)
  wire [49:0] lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2414" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3960" *)
  wire [7:0] lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1645" *)
  reg [7:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2090" *)
  wire [34:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2637" *)
  wire lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4029" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246" *)
  wire [247:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1647" *)
  reg lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1055" *)
  wire [9:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2091" *)
  wire [255:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1633" *)
  reg [7:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2088" *)
  wire [34:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4027" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246" *)
  wire [247:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1634" *)
  reg lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1057" *)
  wire [9:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2089" *)
  wire [255:0] lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1629" *)
  reg [22:0] lut_lookup_3_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3903" *)
  wire [22:0] lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1528" *)
  reg lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1070" *)
  wire lut_lookup_3_FpMantRNE_49U_24U_2_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1641" *)
  reg [22:0] lut_lookup_3_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3900" *)
  wire [22:0] lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1072" *)
  wire lut_lookup_3_FpMantRNE_49U_24U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4107" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4109" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] lut_lookup_3_FpNormalize_8U_49U_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2976" *)
  wire [7:0] lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2138" *)
  wire [48:0] lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2412" *)
  wire [7:0] lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2136" *)
  wire [48:0] lut_lookup_3_FpNormalize_8U_49U_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3590" *)
  wire [30:0] lut_lookup_3_IntLog2_32U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3589" *)
  wire [30:0] lut_lookup_3_IntLog2_32U_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1625" *)
  reg [1:0] lut_lookup_3_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2122" *)
  wire [30:0] lut_lookup_3_IntLog2_32U_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2139" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126" *)
  wire [286:0] lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4062" *)
  wire lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1071" *)
  wire [8:0] lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2137" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126" *)
  wire [286:0] lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4060" *)
  wire lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1540" *)
  reg lut_lookup_3_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2614" *)
  wire lut_lookup_3_else_1_acc_itm_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3883" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_3_else_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1648" *)
  reg [31:0] lut_lookup_3_else_1_else_else_lo_data_f_and_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2107" *)
  wire [34:0] lut_lookup_3_else_1_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1650" *)
  reg lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1651" *)
  reg lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1723" *)
  reg lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1649" *)
  reg lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1785" *)
  wire lut_lookup_3_else_2_and_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1784" *)
  wire lut_lookup_3_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2645" *)
  wire lut_lookup_3_else_else_acc_1_itm_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4077" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_3_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1635" *)
  reg [31:0] lut_lookup_3_else_else_else_else_le_data_f_and_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2106" *)
  wire [34:0] lut_lookup_3_else_else_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2601" *)
  wire lut_lookup_3_else_else_else_if_acc_itm_3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3853" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_3_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2636" *)
  wire lut_lookup_3_else_if_else_if_acc_itm_3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4021" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_3_else_if_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2600" *)
  wire lut_lookup_3_if_else_else_acc_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3851" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] lut_lookup_3_if_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2608" *)
  wire lut_lookup_3_if_else_else_else_else_acc_itm_32_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3867" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_3_if_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3599" *)
  wire [6:0] lut_lookup_3_if_else_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2105" *)
  wire [34:0] lut_lookup_3_if_else_else_else_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3601" *)
  wire [3:0] lut_lookup_3_if_else_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2104" *)
  wire [34:0] lut_lookup_3_if_else_else_else_else_if_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1715" *)
  reg lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1626" *)
  reg [5:0] lut_lookup_3_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2609" *)
  wire lut_lookup_3_if_else_else_else_if_acc_itm_3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3869" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_3_if_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1273" *)
  reg lut_lookup_3_if_else_slc_32_svs_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1274" *)
  reg lut_lookup_3_if_else_slc_32_svs_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1275" *)
  reg lut_lookup_3_if_else_slc_32_svs_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1276" *)
  reg lut_lookup_3_if_else_slc_32_svs_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1713" *)
  reg lut_lookup_3_if_else_slc_32_svs_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2630" *)
  wire lut_lookup_3_if_if_else_acc_itm_9_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3995" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8" *)
  wire [9:0] lut_lookup_3_if_if_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2642" *)
  wire lut_lookup_3_if_if_else_else_if_acc_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4071" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_3_if_if_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1655" *)
  reg lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1656" *)
  reg lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2819" *)
  wire [49:0] lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2821" *)
  wire [49:0] lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2659" *)
  wire lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4121" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2663" *)
  wire lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4129" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1029" *)
  wire lut_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1668" *)
  reg lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1669" *)
  reg lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4593" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4582" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2829" *)
  wire [49:0] lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2827" *)
  wire [49:0] lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2623" *)
  wire lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3925" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3028" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2627" *)
  wire lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3982" *)
  (* unused_bits = "0 1 2 3 4 5 6" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3985" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1027" *)
  wire lut_lookup_4_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2207" *)
  wire lut_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2391" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2389" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2823" *)
  wire [49:0] lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2825" *)
  wire [49:0] lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2407" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3976" *)
  wire [7:0] lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1676" *)
  reg [7:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2094" *)
  wire [34:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2639" *)
  wire lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4040" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246" *)
  wire [247:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1678" *)
  reg lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1051" *)
  wire [9:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2095" *)
  wire [255:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1663" *)
  reg [7:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2092" *)
  wire [34:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4038" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246" *)
  wire [247:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1664" *)
  reg lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1053" *)
  wire [9:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2093" *)
  wire [255:0] lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1659" *)
  reg [22:0] lut_lookup_4_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3909" *)
  wire [22:0] lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1558" *)
  reg lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1067" *)
  wire lut_lookup_4_FpMantRNE_49U_24U_2_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1672" *)
  reg [22:0] lut_lookup_4_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3906" *)
  wire [22:0] lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1069" *)
  wire lut_lookup_4_FpMantRNE_49U_24U_else_and_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4111" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4113" *)
  (* unused_bits = "0 1 2 3 4 5 6 7" *)
  wire [8:0] lut_lookup_4_FpNormalize_8U_49U_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3026" *)
  wire [7:0] lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2142" *)
  wire [48:0] lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2405" *)
  wire [7:0] lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2140" *)
  wire [48:0] lut_lookup_4_FpNormalize_8U_49U_else_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3651" *)
  wire [30:0] lut_lookup_4_IntLog2_32U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3650" *)
  wire [30:0] lut_lookup_4_IntLog2_32U_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1653" *)
  reg [1:0] lut_lookup_4_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2125" *)
  wire [30:0] lut_lookup_4_IntLog2_32U_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2143" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126" *)
  wire [286:0] lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4066" *)
  wire lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1068" *)
  wire [8:0] lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2141" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126" *)
  wire [286:0] lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4064" *)
  wire lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1570" *)
  reg lut_lookup_4_and_svs_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2615" *)
  wire lut_lookup_4_else_1_acc_itm_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3885" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_4_else_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1679" *)
  reg [31:0] lut_lookup_4_else_1_else_else_lo_data_f_and_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2111" *)
  wire [34:0] lut_lookup_4_else_1_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1681" *)
  reg lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1682" *)
  reg lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1735" *)
  reg lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1680" *)
  reg lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1788" *)
  wire lut_lookup_4_else_2_and_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1787" *)
  wire lut_lookup_4_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2647" *)
  wire lut_lookup_4_else_else_acc_1_itm_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4081" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_4_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1665" *)
  reg [31:0] lut_lookup_4_else_else_else_else_le_data_f_and_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2110" *)
  wire [34:0] lut_lookup_4_else_else_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2603" *)
  wire lut_lookup_4_else_else_else_if_acc_itm_3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3857" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_4_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2638" *)
  wire lut_lookup_4_else_if_else_if_acc_itm_3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4032" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_4_else_if_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2602" *)
  wire lut_lookup_4_if_else_else_acc_itm_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3855" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9" *)
  wire [10:0] lut_lookup_4_if_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2610" *)
  wire lut_lookup_4_if_else_else_else_else_acc_itm_32_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3871" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [32:0] lut_lookup_4_if_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3660" *)
  wire [6:0] lut_lookup_4_if_else_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2109" *)
  wire [34:0] lut_lookup_4_if_else_else_else_else_else_rshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3662" *)
  wire [3:0] lut_lookup_4_if_else_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2108" *)
  wire [34:0] lut_lookup_4_if_else_else_else_else_if_lshift_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1728" *)
  reg lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1654" *)
  reg [5:0] lut_lookup_4_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2611" *)
  wire lut_lookup_4_if_else_else_else_if_acc_itm_3_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3873" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_4_if_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1269" *)
  reg lut_lookup_4_if_else_slc_32_svs_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1270" *)
  reg lut_lookup_4_if_else_slc_32_svs_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1271" *)
  reg lut_lookup_4_if_else_slc_32_svs_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1272" *)
  reg lut_lookup_4_if_else_slc_32_svs_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1726" *)
  reg lut_lookup_4_if_else_slc_32_svs_st_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2631" *)
  wire lut_lookup_4_if_if_else_acc_itm_9_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3997" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8" *)
  wire [9:0] lut_lookup_4_if_if_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2643" *)
  wire lut_lookup_4_if_if_else_else_if_acc_itm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4073" *)
  (* unused_bits = "0 1 2" *)
  wire [3:0] lut_lookup_4_if_if_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2477" *)
  wire lut_lookup_FpAdd_8U_23U_1_or_11_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2479" *)
  wire lut_lookup_FpAdd_8U_23U_2_or_10_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2482" *)
  wire lut_lookup_FpAdd_8U_23U_2_or_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2480" *)
  wire lut_lookup_FpAdd_8U_23U_2_or_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2036" *)
  wire lut_lookup_and_112_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2037" *)
  wire lut_lookup_and_113_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2029" *)
  wire lut_lookup_and_118_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2030" *)
  wire lut_lookup_and_119_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2026" *)
  wire lut_lookup_and_120_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2027" *)
  wire lut_lookup_and_121_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2022" *)
  wire lut_lookup_and_122_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2023" *)
  wire lut_lookup_and_123_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2019" *)
  wire lut_lookup_and_124_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2020" *)
  wire lut_lookup_and_125_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2015" *)
  wire lut_lookup_and_126_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2016" *)
  wire lut_lookup_and_127_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1889" *)
  wire lut_lookup_and_132_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1890" *)
  wire lut_lookup_and_133_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1887" *)
  wire lut_lookup_and_134_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1888" *)
  wire lut_lookup_and_135_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1885" *)
  wire lut_lookup_and_136_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1886" *)
  wire lut_lookup_and_137_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1883" *)
  wire lut_lookup_and_138_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1884" *)
  wire lut_lookup_and_139_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2274" *)
  wire lut_lookup_and_13_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2275" *)
  wire lut_lookup_and_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2276" *)
  wire lut_lookup_and_15_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2278" *)
  wire lut_lookup_and_21_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2279" *)
  wire lut_lookup_and_22_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2280" *)
  wire lut_lookup_and_23_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2282" *)
  wire lut_lookup_and_29_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2283" *)
  wire lut_lookup_and_30_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2284" *)
  wire lut_lookup_and_31_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2270" *)
  wire lut_lookup_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2271" *)
  wire lut_lookup_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2272" *)
  wire lut_lookup_and_7_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2574" *)
  wire lut_lookup_else_1_and_13_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2556" *)
  wire lut_lookup_else_1_and_16_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2591" *)
  wire lut_lookup_else_1_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2582" *)
  wire lut_lookup_else_1_and_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2116" *)
  wire [8:0] lut_lookup_else_1_else_else_mux1h_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1475" *)
  reg [31:0] lut_lookup_else_1_lo_index_u_1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1477" *)
  reg [31:0] lut_lookup_else_1_lo_index_u_1_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1505" *)
  reg [31:0] lut_lookup_else_1_lo_index_u_2_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1507" *)
  reg [31:0] lut_lookup_else_1_lo_index_u_2_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1535" *)
  reg [31:0] lut_lookup_else_1_lo_index_u_3_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1537" *)
  reg [31:0] lut_lookup_else_1_lo_index_u_3_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1565" *)
  reg [31:0] lut_lookup_else_1_lo_index_u_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1567" *)
  reg [31:0] lut_lookup_else_1_lo_index_u_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1683" *)
  reg lut_lookup_else_1_lut_lookup_else_1_and_10_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1598" *)
  reg lut_lookup_else_1_lut_lookup_else_1_and_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1624" *)
  reg lut_lookup_else_1_lut_lookup_else_1_and_4_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1652" *)
  reg lut_lookup_else_1_lut_lookup_else_1_and_7_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2486" *)
  wire lut_lookup_else_1_lut_lookup_lo_uflow_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1388" *)
  reg lut_lookup_else_1_slc_32_mdf_1_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1389" *)
  reg lut_lookup_else_1_slc_32_mdf_1_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1390" *)
  reg lut_lookup_else_1_slc_32_mdf_1_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1391" *)
  reg lut_lookup_else_1_slc_32_mdf_1_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1356" *)
  reg lut_lookup_else_1_slc_32_mdf_2_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1357" *)
  reg lut_lookup_else_1_slc_32_mdf_2_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1358" *)
  reg lut_lookup_else_1_slc_32_mdf_2_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1359" *)
  reg lut_lookup_else_1_slc_32_mdf_2_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1324" *)
  reg lut_lookup_else_1_slc_32_mdf_3_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1325" *)
  reg lut_lookup_else_1_slc_32_mdf_3_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1326" *)
  reg lut_lookup_else_1_slc_32_mdf_3_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1327" *)
  reg lut_lookup_else_1_slc_32_mdf_3_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1292" *)
  reg lut_lookup_else_1_slc_32_mdf_sva_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1293" *)
  reg lut_lookup_else_1_slc_32_mdf_sva_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1294" *)
  reg lut_lookup_else_1_slc_32_mdf_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1295" *)
  reg lut_lookup_else_1_slc_32_mdf_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4203" *)
  wire lut_lookup_else_2_else_else_else_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4210" *)
  wire lut_lookup_else_2_else_else_else_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4217" *)
  wire lut_lookup_else_2_else_else_else_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4224" *)
  wire lut_lookup_else_2_else_else_else_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2760" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2754" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1789" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2777" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2771" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1801" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2726" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2720" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1797" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2743" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2737" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1793" *)
  wire lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1686" *)
  reg lut_lookup_else_2_else_else_if_mux_12_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2199" *)
  wire lut_lookup_else_2_else_else_if_mux_12_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1685" *)
  reg lut_lookup_else_2_else_else_if_mux_19_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2200" *)
  wire lut_lookup_else_2_else_else_if_mux_19_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1684" *)
  reg lut_lookup_else_2_else_else_if_mux_26_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2201" *)
  wire lut_lookup_else_2_else_else_if_mux_26_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1687" *)
  reg lut_lookup_else_2_else_else_if_mux_5_itm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2198" *)
  wire lut_lookup_else_2_else_else_if_mux_5_itm_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2725" *)
  wire lut_lookup_else_2_else_else_mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2719" *)
  wire lut_lookup_else_2_else_else_mux_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2714" *)
  wire lut_lookup_else_2_else_else_mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2704" *)
  wire lut_lookup_else_2_else_else_mux_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2742" *)
  wire lut_lookup_else_2_else_else_mux_26_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2736" *)
  wire lut_lookup_else_2_else_else_mux_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2731" *)
  wire lut_lookup_else_2_else_else_mux_28_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2707" *)
  wire lut_lookup_else_2_else_else_mux_33_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2701" *)
  wire lut_lookup_else_2_else_else_mux_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2759" *)
  wire lut_lookup_else_2_else_else_mux_41_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2753" *)
  wire lut_lookup_else_2_else_else_mux_42_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2748" *)
  wire lut_lookup_else_2_else_else_mux_43_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2710" *)
  wire lut_lookup_else_2_else_else_mux_48_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2776" *)
  wire lut_lookup_else_2_else_else_mux_56_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2770" *)
  wire lut_lookup_else_2_else_else_mux_57_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2765" *)
  wire lut_lookup_else_2_else_else_mux_58_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2690" *)
  wire lut_lookup_else_2_else_else_mux_59_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2686" *)
  wire lut_lookup_else_2_else_else_mux_60_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2682" *)
  wire lut_lookup_else_2_else_else_mux_61_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2694" *)
  wire lut_lookup_else_2_else_else_mux_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2242" *)
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2248" *)
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2249" *)
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2255" *)
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2256" *)
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2262" *)
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2263" *)
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_7_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2243" *)
  wire lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2257" *)
  wire lut_lookup_else_2_else_if_mux_12_cse_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2264" *)
  wire lut_lookup_else_2_else_if_mux_17_cse_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2241" *)
  wire lut_lookup_else_2_else_if_mux_2_cse_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2250" *)
  wire lut_lookup_else_2_else_if_mux_7_cse_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2685" *)
  wire lut_lookup_else_2_else_lut_lookup_else_2_else_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2689" *)
  wire lut_lookup_else_2_else_lut_lookup_else_2_else_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2693" *)
  wire lut_lookup_else_2_else_lut_lookup_else_2_else_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2681" *)
  wire lut_lookup_else_2_else_lut_lookup_else_2_else_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2724" *)
  wire lut_lookup_else_2_else_mux_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2718" *)
  wire lut_lookup_else_2_else_mux_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2713" *)
  wire lut_lookup_else_2_else_mux_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2703" *)
  wire lut_lookup_else_2_else_mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2741" *)
  wire lut_lookup_else_2_else_mux_36_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2735" *)
  wire lut_lookup_else_2_else_mux_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2730" *)
  wire lut_lookup_else_2_else_mux_38_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2700" *)
  wire lut_lookup_else_2_else_mux_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2706" *)
  wire lut_lookup_else_2_else_mux_43_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2758" *)
  wire lut_lookup_else_2_else_mux_56_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2752" *)
  wire lut_lookup_else_2_else_mux_57_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2747" *)
  wire lut_lookup_else_2_else_mux_58_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2709" *)
  wire lut_lookup_else_2_else_mux_63_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2775" *)
  wire lut_lookup_else_2_else_mux_76_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2769" *)
  wire lut_lookup_else_2_else_mux_77_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2764" *)
  wire lut_lookup_else_2_else_mux_78_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2717" *)
  wire lut_lookup_else_2_if_lut_lookup_else_2_if_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2740" *)
  wire lut_lookup_else_2_if_lut_lookup_else_2_if_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2734" *)
  wire lut_lookup_else_2_if_lut_lookup_else_2_if_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2757" *)
  wire lut_lookup_else_2_if_lut_lookup_else_2_if_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2751" *)
  wire lut_lookup_else_2_if_lut_lookup_else_2_if_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2774" *)
  wire lut_lookup_else_2_if_lut_lookup_else_2_if_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2768" *)
  wire lut_lookup_else_2_if_lut_lookup_else_2_if_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2723" *)
  wire lut_lookup_else_2_if_lut_lookup_else_2_if_and_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2684" *)
  wire lut_lookup_else_2_if_mux_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2688" *)
  wire lut_lookup_else_2_if_mux_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2692" *)
  wire lut_lookup_else_2_if_mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4202" *)
  wire lut_lookup_else_2_if_mux_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4209" *)
  wire lut_lookup_else_2_if_mux_32_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4216" *)
  wire lut_lookup_else_2_if_mux_33_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4223" *)
  wire lut_lookup_else_2_if_mux_34_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2680" *)
  wire lut_lookup_else_2_if_mux_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2695" *)
  wire lut_lookup_else_2_lut_lookup_else_2_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2696" *)
  wire lut_lookup_else_2_lut_lookup_else_2_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2697" *)
  wire lut_lookup_else_2_lut_lookup_else_2_and_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2698" *)
  wire lut_lookup_else_2_lut_lookup_else_2_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2699" *)
  wire lut_lookup_else_2_mux_103_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2702" *)
  wire lut_lookup_else_2_mux_104_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2705" *)
  wire lut_lookup_else_2_mux_105_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2708" *)
  wire lut_lookup_else_2_mux_106_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2712" *)
  wire lut_lookup_else_2_mux_107_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2716" *)
  wire lut_lookup_else_2_mux_108_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2722" *)
  wire lut_lookup_else_2_mux_109_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2729" *)
  wire lut_lookup_else_2_mux_110_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2733" *)
  wire lut_lookup_else_2_mux_111_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2739" *)
  wire lut_lookup_else_2_mux_112_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2746" *)
  wire lut_lookup_else_2_mux_113_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2750" *)
  wire lut_lookup_else_2_mux_114_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2756" *)
  wire lut_lookup_else_2_mux_115_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2763" *)
  wire lut_lookup_else_2_mux_116_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2767" *)
  wire lut_lookup_else_2_mux_117_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2773" *)
  wire lut_lookup_else_2_mux_118_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2679" *)
  wire lut_lookup_else_2_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2683" *)
  wire lut_lookup_else_2_mux_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2687" *)
  wire lut_lookup_else_2_mux_53_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2691" *)
  wire lut_lookup_else_2_mux_79_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2519" *)
  wire lut_lookup_else_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2579" *)
  wire lut_lookup_else_else_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2581" *)
  wire lut_lookup_else_else_and_9_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2577" *)
  wire lut_lookup_else_else_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1400" *)
  reg lut_lookup_else_else_else_asn_mdf_1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1401" *)
  reg lut_lookup_else_else_else_asn_mdf_1_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1696" *)
  reg lut_lookup_else_else_else_asn_mdf_1_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1368" *)
  reg lut_lookup_else_else_else_asn_mdf_2_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1369" *)
  reg lut_lookup_else_else_else_asn_mdf_2_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1708" *)
  reg lut_lookup_else_else_else_asn_mdf_2_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1336" *)
  reg lut_lookup_else_else_else_asn_mdf_3_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1337" *)
  reg lut_lookup_else_else_else_asn_mdf_3_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1718" *)
  reg lut_lookup_else_else_else_asn_mdf_3_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1304" *)
  reg lut_lookup_else_else_else_asn_mdf_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1305" *)
  reg lut_lookup_else_else_else_asn_mdf_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1731" *)
  reg lut_lookup_else_else_else_asn_mdf_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1910" *)
  wire [8:0] lut_lookup_else_else_else_else_mux1h_1_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1912" *)
  wire [8:0] lut_lookup_else_else_else_else_mux1h_2_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1914" *)
  wire [8:0] lut_lookup_else_else_else_else_mux1h_3_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1908" *)
  wire [8:0] lut_lookup_else_else_else_else_mux1h_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1458" *)
  reg [31:0] lut_lookup_else_else_else_le_index_u_1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1459" *)
  reg [31:0] lut_lookup_else_else_else_le_index_u_1_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1489" *)
  reg [31:0] lut_lookup_else_else_else_le_index_u_2_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1490" *)
  reg [31:0] lut_lookup_else_else_else_le_index_u_2_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1519" *)
  reg [31:0] lut_lookup_else_else_else_le_index_u_3_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1520" *)
  reg [31:0] lut_lookup_else_else_else_le_index_u_3_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1549" *)
  reg [31:0] lut_lookup_else_else_else_le_index_u_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1550" *)
  reg [31:0] lut_lookup_else_else_else_le_index_u_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3777" *)
  wire [5:0] lut_lookup_else_else_else_lut_lookup_else_else_else_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3789" *)
  wire [5:0] lut_lookup_else_else_else_lut_lookup_else_else_else_and_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3800" *)
  wire [5:0] lut_lookup_else_else_else_lut_lookup_else_else_else_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3811" *)
  wire [5:0] lut_lookup_else_else_else_lut_lookup_else_else_else_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1667" *)
  reg lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3249" *)
  wire lut_lookup_else_else_lut_lookup_else_else_and_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1585" *)
  reg lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3259" *)
  wire lut_lookup_else_else_lut_lookup_else_else_and_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1611" *)
  reg lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3256" *)
  wire lut_lookup_else_else_lut_lookup_else_else_and_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1637" *)
  reg lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3252" *)
  wire lut_lookup_else_else_lut_lookup_else_else_and_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2470" *)
  wire lut_lookup_else_else_lut_lookup_else_else_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1402" *)
  reg lut_lookup_else_else_slc_32_mdf_1_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1403" *)
  reg lut_lookup_else_else_slc_32_mdf_1_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1370" *)
  reg lut_lookup_else_else_slc_32_mdf_2_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1371" *)
  reg lut_lookup_else_else_slc_32_mdf_2_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1338" *)
  reg lut_lookup_else_else_slc_32_mdf_3_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1339" *)
  reg lut_lookup_else_else_slc_32_mdf_3_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1306" *)
  reg lut_lookup_else_else_slc_32_mdf_sva_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1307" *)
  reg lut_lookup_else_else_slc_32_mdf_sva_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1404" *)
  reg [34:0] lut_lookup_else_if_else_le_fra_1_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1372" *)
  reg [34:0] lut_lookup_else_if_else_le_fra_2_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1340" *)
  reg [34:0] lut_lookup_else_if_else_le_fra_3_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1308" *)
  reg [34:0] lut_lookup_else_if_else_le_fra_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1817" *)
  wire [8:0] lut_lookup_else_if_else_le_int_1_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1816" *)
  wire [8:0] lut_lookup_else_if_else_le_int_2_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1815" *)
  wire [8:0] lut_lookup_else_if_else_le_int_3_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1814" *)
  wire [8:0] lut_lookup_else_if_else_le_int_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1309" *)
  reg lut_lookup_else_if_lor_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1310" *)
  reg lut_lookup_else_if_lor_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2195" *)
  wire lut_lookup_else_if_lor_1_lpi_1_dfm_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1730" *)
  reg lut_lookup_else_if_lor_1_lpi_1_dfm_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1405" *)
  reg lut_lookup_else_if_lor_5_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1406" *)
  reg lut_lookup_else_if_lor_5_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1906" *)
  wire lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1695" *)
  reg lut_lookup_else_if_lor_5_lpi_1_dfm_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1373" *)
  reg lut_lookup_else_if_lor_6_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1374" *)
  reg lut_lookup_else_if_lor_6_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2191" *)
  wire lut_lookup_else_if_lor_6_lpi_1_dfm_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1707" *)
  reg lut_lookup_else_if_lor_6_lpi_1_dfm_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1341" *)
  reg lut_lookup_else_if_lor_7_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1342" *)
  reg lut_lookup_else_if_lor_7_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2193" *)
  wire lut_lookup_else_if_lor_7_lpi_1_dfm_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1717" *)
  reg lut_lookup_else_if_lor_7_lpi_1_dfm_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2762" *)
  wire [5:0] lut_lookup_else_if_lut_lookup_else_if_and_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2711" *)
  wire [5:0] lut_lookup_else_if_lut_lookup_else_if_and_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2728" *)
  wire [5:0] lut_lookup_else_if_lut_lookup_else_if_and_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2745" *)
  wire [5:0] lut_lookup_else_if_lut_lookup_else_if_and_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4013" *)
  wire lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4024" *)
  wire lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4036" *)
  wire lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4002" *)
  wire lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2594" *)
  wire lut_lookup_else_if_oelse_1_and_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2595" *)
  wire lut_lookup_else_if_oelse_1_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2588" *)
  wire lut_lookup_else_if_oelse_1_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1666" *)
  reg lut_lookup_else_mux_129_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4001" *)
  wire lut_lookup_else_mux_172_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4012" *)
  wire lut_lookup_else_mux_174_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4023" *)
  wire lut_lookup_else_mux_176_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4035" *)
  wire lut_lookup_else_mux_178_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1858" *)
  wire lut_lookup_else_mux_180_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1859" *)
  wire lut_lookup_else_mux_182_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1860" *)
  wire lut_lookup_else_mux_184_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1861" *)
  wire lut_lookup_else_mux_186_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1610" *)
  reg lut_lookup_else_mux_43_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1636" *)
  reg lut_lookup_else_mux_86_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1584" *)
  reg lut_lookup_else_mux_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1285" *)
  reg lut_lookup_else_unequal_tmp_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1286" *)
  reg lut_lookup_else_unequal_tmp_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1287" *)
  reg lut_lookup_else_unequal_tmp_18;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1392" *)
  reg [34:0] lut_lookup_if_1_else_lo_fra_1_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1360" *)
  reg [34:0] lut_lookup_if_1_else_lo_fra_2_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1328" *)
  reg [34:0] lut_lookup_if_1_else_lo_fra_3_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1296" *)
  reg [34:0] lut_lookup_if_1_else_lo_fra_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2245" *)
  wire [8:0] lut_lookup_if_1_else_lo_int_1_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2252" *)
  wire [8:0] lut_lookup_if_1_else_lo_int_2_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2259" *)
  wire [8:0] lut_lookup_if_1_else_lo_int_3_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2266" *)
  wire [8:0] lut_lookup_if_1_else_lo_int_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1297" *)
  reg lut_lookup_if_1_lor_1_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1298" *)
  reg lut_lookup_if_1_lor_1_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2196" *)
  wire lut_lookup_if_1_lor_1_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1734" *)
  reg lut_lookup_if_1_lor_1_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1393" *)
  reg lut_lookup_if_1_lor_5_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1394" *)
  reg lut_lookup_if_1_lor_5_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1700" *)
  reg lut_lookup_if_1_lor_5_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1361" *)
  reg lut_lookup_if_1_lor_6_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1362" *)
  reg lut_lookup_if_1_lor_6_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2192" *)
  wire lut_lookup_if_1_lor_6_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1711" *)
  reg lut_lookup_if_1_lor_6_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1329" *)
  reg lut_lookup_if_1_lor_7_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1330" *)
  reg lut_lookup_if_1_lor_7_lpi_1_dfm_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2194" *)
  wire lut_lookup_if_1_lor_7_lpi_1_dfm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1722" *)
  reg lut_lookup_if_1_lor_7_lpi_1_dfm_st_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4003" *)
  wire lut_lookup_if_1_lut_lookup_if_1_and_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4014" *)
  wire lut_lookup_if_1_lut_lookup_if_1_and_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4025" *)
  wire lut_lookup_if_1_lut_lookup_if_1_and_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4034" *)
  wire lut_lookup_if_1_lut_lookup_if_1_and_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2578" *)
  wire lut_lookup_if_1_oelse_1_and_12_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2589" *)
  wire lut_lookup_if_1_oelse_1_and_14_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2586" *)
  wire lut_lookup_if_1_oelse_1_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2587" *)
  wire lut_lookup_if_1_oelse_1_and_5_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2593" *)
  wire lut_lookup_if_1_oelse_1_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2738" *)
  wire lut_lookup_if_2_lut_lookup_if_2_and_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2744" *)
  wire lut_lookup_if_2_lut_lookup_if_2_and_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2755" *)
  wire lut_lookup_if_2_lut_lookup_if_2_and_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2761" *)
  wire lut_lookup_if_2_lut_lookup_if_2_and_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2772" *)
  wire lut_lookup_if_2_lut_lookup_if_2_and_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2778" *)
  wire lut_lookup_if_2_lut_lookup_if_2_and_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2721" *)
  wire lut_lookup_if_2_lut_lookup_if_2_and_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2727" *)
  wire lut_lookup_if_2_lut_lookup_if_2_and_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2715" *)
  wire lut_lookup_if_2_mux_21_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2732" *)
  wire lut_lookup_if_2_mux_22_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2749" *)
  wire lut_lookup_if_2_mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2766" *)
  wire lut_lookup_if_2_mux_24_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1412" *)
  reg lut_lookup_if_else_else_else_asn_mdf_1_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1380" *)
  reg lut_lookup_if_else_else_else_asn_mdf_2_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1348" *)
  reg lut_lookup_if_else_else_else_asn_mdf_3_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1316" *)
  reg lut_lookup_if_else_else_else_asn_mdf_sva_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2561" *)
  wire lut_lookup_if_else_else_else_else_if_lut_lookup_if_else_else_else_else_if_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3240" *)
  wire [34:0] lut_lookup_if_else_else_else_else_mux_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3241" *)
  wire [34:0] lut_lookup_if_else_else_else_else_mux_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3242" *)
  wire [34:0] lut_lookup_if_else_else_else_else_mux_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3239" *)
  wire [34:0] lut_lookup_if_else_else_else_else_mux_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1951" *)
  wire [8:0] lut_lookup_if_else_else_else_le_index_s_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1953" *)
  wire [8:0] lut_lookup_if_else_else_else_le_index_s_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1955" *)
  wire [8:0] lut_lookup_if_else_else_else_le_index_s_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1957" *)
  wire [8:0] lut_lookup_if_else_else_else_le_index_s_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1744" *)
  reg [30:0] lut_lookup_if_else_else_le_data_sub_1_sva_1_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2210" *)
  wire [31:0] lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1745" *)
  reg [30:0] lut_lookup_if_else_else_le_data_sub_2_sva_1_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2212" *)
  wire [31:0] lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1746" *)
  reg [30:0] lut_lookup_if_else_else_le_data_sub_3_sva_1_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2214" *)
  wire [31:0] lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1747" *)
  reg [30:0] lut_lookup_if_else_else_le_data_sub_sva_1_30_0_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2216" *)
  wire [31:0] lut_lookup_if_else_else_le_data_sub_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1413" *)
  reg lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1414" *)
  reg lut_lookup_if_else_else_slc_10_mdf_1_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1691" *)
  reg lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1381" *)
  reg lut_lookup_if_else_else_slc_10_mdf_2_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1382" *)
  reg lut_lookup_if_else_else_slc_10_mdf_2_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1703" *)
  reg lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1349" *)
  reg lut_lookup_if_else_else_slc_10_mdf_3_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1350" *)
  reg lut_lookup_if_else_else_slc_10_mdf_3_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1714" *)
  reg lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1317" *)
  reg lut_lookup_if_else_else_slc_10_mdf_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1318" *)
  reg lut_lookup_if_else_else_slc_10_mdf_sva_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1727" *)
  reg lut_lookup_if_else_else_slc_10_mdf_sva_st_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2570" *)
  wire lut_lookup_if_else_if_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2562" *)
  wire lut_lookup_if_else_if_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3250" *)
  wire lut_lookup_if_else_lut_lookup_if_else_and_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3253" *)
  wire lut_lookup_if_else_lut_lookup_if_else_and_12_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3257" *)
  wire lut_lookup_if_else_lut_lookup_if_else_and_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3260" *)
  wire lut_lookup_if_else_lut_lookup_if_else_and_14_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1897" *)
  wire lut_lookup_if_else_lut_lookup_if_else_or_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1898" *)
  wire lut_lookup_if_else_lut_lookup_if_else_or_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1899" *)
  wire lut_lookup_if_else_lut_lookup_if_else_or_3_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1896" *)
  wire lut_lookup_if_else_lut_lookup_if_else_or_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1824" *)
  wire [8:0] lut_lookup_if_if_else_else_le_index_s_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1822" *)
  wire [8:0] lut_lookup_if_if_else_else_le_index_s_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1820" *)
  wire [8:0] lut_lookup_if_if_else_else_le_index_s_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1818" *)
  wire [8:0] lut_lookup_if_if_else_else_le_index_s_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1244" *)
  reg lut_lookup_if_if_lor_1_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2218" *)
  wire lut_lookup_if_if_lor_1_lpi_1_dfm_mx0w3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1264" *)
  reg lut_lookup_if_if_lor_5_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2222" *)
  wire lut_lookup_if_if_lor_5_lpi_1_dfm_mx0w3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1257" *)
  reg lut_lookup_if_if_lor_6_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2221" *)
  wire lut_lookup_if_if_lor_6_lpi_1_dfm_mx0w3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1251" *)
  reg lut_lookup_if_if_lor_7_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2220" *)
  wire lut_lookup_if_if_lor_7_lpi_1_dfm_mx0w3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3251" *)
  wire lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3254" *)
  wire lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3258" *)
  wire lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3261" *)
  wire lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3877" *)
  wire lut_lookup_if_if_lut_lookup_if_if_or_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3876" *)
  wire lut_lookup_if_if_lut_lookup_if_if_or_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3875" *)
  wire lut_lookup_if_if_lut_lookup_if_if_or_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3878" *)
  wire lut_lookup_if_if_lut_lookup_if_if_or_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2569" *)
  wire lut_lookup_if_if_oelse_1_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1810" *)
  wire lut_lookup_if_mux_123_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1812" *)
  wire lut_lookup_if_mux_41_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1811" *)
  wire lut_lookup_if_mux_82_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1813" *)
  wire lut_lookup_if_mux_mx0w1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2202" *)
  wire lut_lookup_if_unequal_tmp_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1739" *)
  reg [22:0] lut_lookup_le_fraction_1_lpi_1_dfm_16_34_12_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1399" *)
  reg [34:0] lut_lookup_le_fraction_1_lpi_1_dfm_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1411" *)
  reg [34:0] lut_lookup_le_fraction_1_lpi_1_dfm_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2244" *)
  wire [34:0] lut_lookup_le_fraction_1_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1738" *)
  reg [22:0] lut_lookup_le_fraction_2_lpi_1_dfm_16_34_12_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1367" *)
  reg [34:0] lut_lookup_le_fraction_2_lpi_1_dfm_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1379" *)
  reg [34:0] lut_lookup_le_fraction_2_lpi_1_dfm_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2251" *)
  wire [34:0] lut_lookup_le_fraction_2_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1737" *)
  reg [22:0] lut_lookup_le_fraction_3_lpi_1_dfm_16_34_12_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1335" *)
  reg [34:0] lut_lookup_le_fraction_3_lpi_1_dfm_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1347" *)
  reg [34:0] lut_lookup_le_fraction_3_lpi_1_dfm_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2258" *)
  wire [34:0] lut_lookup_le_fraction_3_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1736" *)
  reg [22:0] lut_lookup_le_fraction_lpi_1_dfm_16_34_12_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1303" *)
  reg [34:0] lut_lookup_le_fraction_lpi_1_dfm_21;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1315" *)
  reg [34:0] lut_lookup_le_fraction_lpi_1_dfm_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2265" *)
  wire [34:0] lut_lookup_le_fraction_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1397" *)
  reg [5:0] lut_lookup_le_index_0_5_0_1_lpi_1_dfm_25;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1398" *)
  reg [5:0] lut_lookup_le_index_0_5_0_1_lpi_1_dfm_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1409" *)
  reg [5:0] lut_lookup_le_index_0_5_0_1_lpi_1_dfm_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1410" *)
  reg [5:0] lut_lookup_le_index_0_5_0_1_lpi_1_dfm_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1415" *)
  reg [5:0] lut_lookup_le_index_0_5_0_1_lpi_1_dfm_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1365" *)
  reg [5:0] lut_lookup_le_index_0_5_0_2_lpi_1_dfm_25;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1366" *)
  reg [5:0] lut_lookup_le_index_0_5_0_2_lpi_1_dfm_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1377" *)
  reg [5:0] lut_lookup_le_index_0_5_0_2_lpi_1_dfm_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1378" *)
  reg [5:0] lut_lookup_le_index_0_5_0_2_lpi_1_dfm_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1383" *)
  reg [5:0] lut_lookup_le_index_0_5_0_2_lpi_1_dfm_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1333" *)
  reg [5:0] lut_lookup_le_index_0_5_0_3_lpi_1_dfm_25;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1334" *)
  reg [5:0] lut_lookup_le_index_0_5_0_3_lpi_1_dfm_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1345" *)
  reg [5:0] lut_lookup_le_index_0_5_0_3_lpi_1_dfm_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1346" *)
  reg [5:0] lut_lookup_le_index_0_5_0_3_lpi_1_dfm_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1351" *)
  reg [5:0] lut_lookup_le_index_0_5_0_3_lpi_1_dfm_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1301" *)
  reg [5:0] lut_lookup_le_index_0_5_0_lpi_1_dfm_25;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1302" *)
  reg [5:0] lut_lookup_le_index_0_5_0_lpi_1_dfm_26;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1313" *)
  reg [5:0] lut_lookup_le_index_0_5_0_lpi_1_dfm_27;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1314" *)
  reg [5:0] lut_lookup_le_index_0_5_0_lpi_1_dfm_28;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1319" *)
  reg [5:0] lut_lookup_le_index_0_5_0_lpi_1_dfm_29;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1803" *)
  wire lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1799" *)
  wire lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1795" *)
  wire lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1791" *)
  wire lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1777" *)
  wire lut_lookup_le_miss_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1780" *)
  wire lut_lookup_le_miss_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1783" *)
  wire lut_lookup_le_miss_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1786" *)
  wire lut_lookup_le_miss_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1460" *)
  reg lut_lookup_le_uflow_1_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1491" *)
  reg lut_lookup_le_uflow_2_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1521" *)
  reg lut_lookup_le_uflow_3_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2469" *)
  wire lut_lookup_le_uflow_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1551" *)
  reg lut_lookup_le_uflow_lpi_1_dfm_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2247" *)
  wire [34:0] lut_lookup_lo_fraction_1_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1387" *)
  reg [34:0] lut_lookup_lo_fraction_1_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2254" *)
  wire [34:0] lut_lookup_lo_fraction_2_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1355" *)
  reg [34:0] lut_lookup_lo_fraction_2_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2261" *)
  wire [34:0] lut_lookup_lo_fraction_3_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1323" *)
  reg [34:0] lut_lookup_lo_fraction_3_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2268" *)
  wire [34:0] lut_lookup_lo_fraction_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1291" *)
  reg [34:0] lut_lookup_lo_fraction_lpi_1_dfm_9;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2246" *)
  wire [7:0] lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1384" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1385" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1386" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2373" *)
  wire [1:0] lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2253" *)
  wire [7:0] lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1352" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1353" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1354" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2374" *)
  wire [1:0] lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2260" *)
  wire [7:0] lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1320" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1321" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1322" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2375" *)
  wire [1:0] lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2267" *)
  wire [7:0] lut_lookup_lo_index_0_7_0_lpi_1_dfm_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1288" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_lpi_1_dfm_11;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1289" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_lpi_1_dfm_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1290" *)
  reg [7:0] lut_lookup_lo_index_0_7_0_lpi_1_dfm_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2376" *)
  wire [1:0] lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1804" *)
  wire lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1800" *)
  wire lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1796" *)
  wire lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1792" *)
  wire lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2471" *)
  wire lut_lookup_lo_index_0_and_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2485" *)
  wire lut_lookup_lo_index_0_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2487" *)
  wire lut_lookup_lo_index_0_and_6_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2488" *)
  wire lut_lookup_lo_index_0_and_8_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2468" *)
  wire lut_lookup_lo_index_0_and_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1802" *)
  wire lut_lookup_lo_miss_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1798" *)
  wire lut_lookup_lo_miss_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1794" *)
  wire lut_lookup_lo_miss_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1790" *)
  wire lut_lookup_lo_miss_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1478" *)
  reg lut_lookup_lo_uflow_1_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1479" *)
  reg lut_lookup_lo_uflow_1_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1508" *)
  reg lut_lookup_lo_uflow_2_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1509" *)
  reg lut_lookup_lo_uflow_2_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1538" *)
  reg lut_lookup_lo_uflow_3_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1539" *)
  reg lut_lookup_lo_uflow_3_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2472" *)
  wire lut_lookup_lo_uflow_and_4_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1568" *)
  reg lut_lookup_lo_uflow_lpi_1_dfm_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1569" *)
  reg lut_lookup_lo_uflow_lpi_1_dfm_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2677" *)
  wire [11:0] lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2675" *)
  wire [11:0] lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2673" *)
  wire [11:0] lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2671" *)
  wire [11:0] lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3476" *)
  wire [22:0] lut_lookup_lut_lookup_mux_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3592" *)
  wire [22:0] lut_lookup_lut_lookup_mux_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3653" *)
  wire [22:0] lut_lookup_lut_lookup_mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3541" *)
  wire [22:0] lut_lookup_lut_lookup_mux_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2281" *)
  wire lut_lookup_lut_lookup_nor_16_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2277" *)
  wire lut_lookup_lut_lookup_nor_17_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2273" *)
  wire lut_lookup_lut_lookup_nor_18_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2269" *)
  wire lut_lookup_lut_lookup_nor_19_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2678" *)
  wire lut_lookup_not_36_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2676" *)
  wire lut_lookup_not_37_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2674" *)
  wire lut_lookup_not_38_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2672" *)
  wire lut_lookup_not_39_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1775" *)
  wire lut_lookup_or_11_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1776" *)
  wire lut_lookup_or_15_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2034" *)
  wire lut_lookup_or_16_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2012" *)
  wire lut_lookup_or_17_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2013" *)
  wire lut_lookup_or_18_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1773" *)
  wire lut_lookup_or_3_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1774" *)
  wire lut_lookup_or_7_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2033" *)
  wire lut_lookup_or_rgt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1461" *)
  reg lut_lookup_unequal_tmp_13;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2219" *)
  wire lut_lookup_unequal_tmp_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1756" *)
  wire main_stage_en_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1237" *)
  reg main_stage_v_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2178" *)
  wire main_stage_v_1_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1238" *)
  reg main_stage_v_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2180" *)
  wire main_stage_v_2_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1239" *)
  reg main_stage_v_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2181" *)
  wire main_stage_v_3_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1240" *)
  reg main_stage_v_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2190" *)
  wire main_stage_v_4_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1241" *)
  reg main_stage_v_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2197" *)
  wire main_stage_v_5_mx0c1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3701" *)
  wire mux_1004_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3703" *)
  wire mux_1013_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3709" *)
  wire mux_1014_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3707" *)
  wire mux_1015_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3713" *)
  wire mux_1031_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3719" *)
  wire mux_1032_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3717" *)
  wire mux_1033_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3723" *)
  wire mux_1049_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3727" *)
  wire mux_1051_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3728" *)
  wire mux_1053_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3729" *)
  wire mux_1055_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3730" *)
  wire mux_1056_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3733" *)
  wire mux_1057_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3731" *)
  wire mux_1058_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3736" *)
  wire mux_1059_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3739" *)
  wire mux_1060_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3742" *)
  wire mux_1061_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3745" *)
  wire mux_1062_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3748" *)
  wire mux_1063_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3751" *)
  wire mux_1064_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3754" *)
  wire mux_1066_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3757" *)
  wire mux_1067_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3762" *)
  wire mux_1068_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3760" *)
  wire mux_1069_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3765" *)
  wire mux_1070_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3768" *)
  wire mux_1071_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3771" *)
  wire mux_1073_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3774" *)
  wire mux_1074_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3779" *)
  wire mux_1075_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3782" *)
  wire mux_1076_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3778" *)
  wire mux_1077_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3785" *)
  wire mux_1078_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3787" *)
  wire mux_1079_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3791" *)
  wire mux_1081_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3794" *)
  wire mux_1083_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3790" *)
  wire mux_1084_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3796" *)
  wire mux_1085_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3798" *)
  wire mux_1086_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3802" *)
  wire mux_1088_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3805" *)
  wire mux_1090_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3801" *)
  wire mux_1091_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3807" *)
  wire mux_1092_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3809" *)
  wire mux_1093_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3813" *)
  wire mux_1094_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3816" *)
  wire mux_1095_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3812" *)
  wire mux_1096_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3819" *)
  wire mux_1097_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3821" *)
  wire mux_1098_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3825" *)
  wire mux_1099_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3824" *)
  wire mux_1100_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3823" *)
  wire mux_1101_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3829" *)
  wire mux_1103_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3830" *)
  wire mux_1104_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3833" *)
  wire mux_1106_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3834" *)
  wire mux_1107_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3837" *)
  wire mux_1110_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3840" *)
  wire mux_1112_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3841" *)
  wire mux_1115_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3842" *)
  wire mux_1118_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2781" *)
  wire mux_1120_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2780" *)
  wire mux_1121_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2532" *)
  wire mux_1122_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2848" *)
  wire mux_1125_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2545" *)
  wire mux_1126_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4161" *)
  wire mux_1129_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3126" *)
  wire mux_1138_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3125" *)
  wire mux_1139_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4171" *)
  wire mux_1140_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4169" *)
  wire mux_1141_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4163" *)
  wire mux_1142_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3156" *)
  wire mux_1151_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3155" *)
  wire mux_1152_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4174" *)
  wire mux_1153_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4172" *)
  wire mux_1154_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4165" *)
  wire mux_1155_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3188" *)
  wire mux_1164_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3187" *)
  wire mux_1165_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4177" *)
  wire mux_1166_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4175" *)
  wire mux_1167_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4167" *)
  wire mux_1168_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3217" *)
  wire mux_1177_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3216" *)
  wire mux_1178_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4180" *)
  wire mux_1179_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4178" *)
  wire mux_1180_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3297" *)
  wire mux_1185_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3321" *)
  wire mux_1186_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2571" *)
  wire mux_1187_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2572" *)
  wire mux_1188_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3496" *)
  wire mux_1189_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3499" *)
  wire mux_1190_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3552" *)
  wire mux_1194_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3555" *)
  wire mux_1195_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3603" *)
  wire mux_1199_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2910" *)
  wire mux_119_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3606" *)
  wire mux_1200_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3664" *)
  wire mux_1204_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3667" *)
  wire mux_1205_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2833" *)
  wire mux_1209_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2912" *)
  wire mux_120_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2835" *)
  wire mux_1210_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2942" *)
  wire mux_1211_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2992" *)
  wire mux_1212_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2838" *)
  wire mux_1218_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2836" *)
  wire mux_1219_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2909" *)
  wire mux_121_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2844" *)
  wire mux_1220_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2852" *)
  wire mux_1222_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2851" *)
  wire mux_1223_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2849" *)
  wire mux_1224_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2896" *)
  wire mux_1225_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2894" *)
  wire mux_1226_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2902" *)
  wire mux_1227_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2907" *)
  wire mux_1229_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2906" *)
  wire mux_1230_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2945" *)
  wire mux_1231_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2943" *)
  wire mux_1232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2952" *)
  wire mux_1233_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4189" *)
  wire mux_1234_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2958" *)
  wire mux_1235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2957" *)
  wire mux_1236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2955" *)
  wire mux_1237_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2995" *)
  wire mux_1238_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2993" *)
  wire mux_1239_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2914" *)
  wire mux_123_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3002" *)
  wire mux_1240_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4192" *)
  wire mux_1241_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3008" *)
  wire mux_1242_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3007" *)
  wire mux_1243_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3005" *)
  wire mux_1244_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3480" *)
  wire mux_1245_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3478" *)
  wire mux_1246_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3519" *)
  wire mux_1247_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3517" *)
  wire mux_1248_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3570" *)
  wire mux_1249_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2919" *)
  wire mux_124_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3569" *)
  wire mux_1250_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3618" *)
  wire mux_1251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3679" *)
  wire mux_1252_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2918" *)
  wire mux_125_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4198" *)
  wire mux_1261_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3693" *)
  wire mux_1266_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3715" *)
  wire mux_1267_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3705" *)
  wire mux_1268_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3670" *)
  wire mux_1269_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2923" *)
  wire mux_126_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3641" *)
  wire mux_1270_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3633" *)
  wire mux_1271_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3609" *)
  wire mux_1278_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3558" *)
  wire mux_1279_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2922" *)
  wire mux_127_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3502" *)
  wire mux_1280_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3465" *)
  wire mux_1281_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3443" *)
  wire mux_1282_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3648" *)
  wire mux_1283_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3629" *)
  wire mux_1284_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2568" *)
  wire mux_1285_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4204" *)
  wire mux_1288_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4205" *)
  wire mux_1289_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2917" *)
  wire mux_128_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4211" *)
  wire mux_1291_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4212" *)
  wire mux_1292_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4218" *)
  wire mux_1294_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4219" *)
  wire mux_1295_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4225" *)
  wire mux_1297_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4226" *)
  wire mux_1298_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2931" *)
  wire mux_130_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2930" *)
  wire mux_131_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2935" *)
  wire mux_132_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2937" *)
  wire mux_133_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2938" *)
  wire mux_134_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2936" *)
  wire mux_135_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2941" *)
  wire mux_137_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2939" *)
  wire mux_138_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2832" *)
  wire mux_13_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2948" *)
  wire mux_141_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2960" *)
  wire mux_155_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2962" *)
  wire mux_156_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2959" *)
  wire mux_157_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2964" *)
  wire mux_159_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2969" *)
  wire mux_160_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2968" *)
  wire mux_161_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2973" *)
  wire mux_162_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2972" *)
  wire mux_163_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2967" *)
  wire mux_164_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2981" *)
  wire mux_165_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2983" *)
  wire mux_166_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2980" *)
  wire mux_167_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2986" *)
  wire mux_169_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2987" *)
  wire mux_170_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2985" *)
  wire mux_171_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2991" *)
  wire mux_173_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2988" *)
  wire mux_174_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2998" *)
  wire mux_177_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4134" *)
  wire mux_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3010" *)
  wire mux_198_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3012" *)
  wire mux_199_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3009" *)
  wire mux_200_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3014" *)
  wire mux_202_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3019" *)
  wire mux_203_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3018" *)
  wire mux_204_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3023" *)
  wire mux_205_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3022" *)
  wire mux_206_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3017" *)
  wire mux_207_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3031" *)
  wire mux_209_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2147" *)
  wire mux_20_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3033" *)
  wire mux_210_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3030" *)
  wire mux_211_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3036" *)
  wire mux_213_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3037" *)
  wire mux_214_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3035" *)
  wire mux_215_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3039" *)
  wire mux_216_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3041" *)
  wire mux_217_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3038" *)
  wire mux_218_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3043" *)
  wire mux_219_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3046" *)
  wire mux_220_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3049" *)
  wire mux_222_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3053" *)
  wire mux_223_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3055" *)
  wire mux_224_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3052" *)
  wire mux_225_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3058" *)
  wire mux_226_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3060" *)
  wire mux_228_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3064" *)
  wire mux_229_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3066" *)
  wire mux_230_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3063" *)
  wire mux_231_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3068" *)
  wire mux_232_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3071" *)
  wire mux_234_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3075" *)
  wire mux_235_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3077" *)
  wire mux_236_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3074" *)
  wire mux_237_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3080" *)
  wire mux_238_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2890" *)
  wire mux_23_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3081" *)
  wire mux_240_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3085" *)
  wire mux_241_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3088" *)
  wire mux_242_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3087" *)
  wire mux_243_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3084" *)
  wire mux_244_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3089" *)
  wire mux_245_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3092" *)
  wire mux_247_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3096" *)
  wire mux_248_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3098" *)
  wire mux_249_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3095" *)
  wire mux_250_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3100" *)
  wire mux_251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3101" *)
  wire mux_253_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3105" *)
  wire mux_254_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3107" *)
  wire mux_255_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3104" *)
  wire mux_256_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3109" *)
  wire mux_257_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3112" *)
  wire mux_259_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2148" *)
  wire mux_25_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3116" *)
  wire mux_260_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3118" *)
  wire mux_261_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3115" *)
  wire mux_262_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3121" *)
  wire mux_263_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3122" *)
  wire mux_265_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3128" *)
  wire mux_267_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3131" *)
  wire mux_268_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3134" *)
  wire mux_269_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2149" *)
  wire mux_26_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3136" *)
  wire mux_270_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3141" *)
  wire mux_272_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3140" *)
  wire mux_273_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3139" *)
  wire mux_274_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3142" *)
  wire mux_275_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3143" *)
  wire mux_276_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3144" *)
  wire mux_277_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3147" *)
  wire mux_278_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3149" *)
  wire mux_279_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2940" *)
  wire mux_27_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3151" *)
  wire mux_281_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2592" *)
  wire mux_283_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3153" *)
  wire mux_284_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3154" *)
  wire mux_285_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3158" *)
  wire mux_286_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3161" *)
  wire mux_287_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3166" *)
  wire mux_288_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3164" *)
  wire mux_289_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3171" *)
  wire mux_290_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3169" *)
  wire mux_291_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4147" *)
  wire mux_292_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3176" *)
  wire mux_294_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3175" *)
  wire mux_295_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3174" *)
  wire mux_296_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3177" *)
  wire mux_297_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3178" *)
  wire mux_299_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4132" *)
  wire mux_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3181" *)
  wire mux_300_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3184" *)
  wire mux_301_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3185" *)
  wire mux_303_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3190" *)
  wire mux_308_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3193" *)
  wire mux_309_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3196" *)
  wire mux_310_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3198" *)
  wire mux_311_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3203" *)
  wire mux_314_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3202" *)
  wire mux_315_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3201" *)
  wire mux_316_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3204" *)
  wire mux_319_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2990" *)
  wire mux_31_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3207" *)
  wire mux_320_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3209" *)
  wire mux_322_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3211" *)
  wire mux_325_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3214" *)
  wire mux_328_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3215" *)
  wire mux_329_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2989" *)
  wire mux_32_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3213" *)
  wire mux_330_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3219" *)
  wire mux_332_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3222" *)
  wire mux_333_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3225" *)
  wire mux_334_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3227" *)
  wire mux_335_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3230" *)
  wire mux_343_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3233" *)
  wire mux_344_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3235" *)
  wire mux_346_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3237" *)
  wire mux_349_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3244" *)
  wire mux_356_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3243" *)
  wire mux_357_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3247" *)
  wire mux_358_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3248" *)
  wire mux_359_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3246" *)
  wire mux_360_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3255" *)
  wire mux_366_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3264" *)
  wire mux_371_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3262" *)
  wire mux_372_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2834" *)
  wire mux_38_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2831" *)
  wire mux_39_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2146" *)
  wire mux_3_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2841" *)
  wire mux_42_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3316" *)
  wire mux_477_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2779" *)
  wire mux_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3329" *)
  wire mux_518_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3335" *)
  wire mux_534_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3343" *)
  wire mux_548_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2854" *)
  wire mux_57_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2528" *)
  wire mux_580_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4148" *)
  wire mux_581_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2150" *)
  wire mux_582_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2856" *)
  wire mux_58_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4149" *)
  wire mux_594_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2151" *)
  wire mux_595_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3301" *)
  wire mux_598_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3300" *)
  wire mux_599_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2853" *)
  wire mux_59_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3299" *)
  wire mux_600_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3305" *)
  wire mux_601_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3304" *)
  wire mux_602_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3303" *)
  wire mux_605_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3298" *)
  wire mux_606_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3310" *)
  wire mux_611_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4153" *)
  wire mux_615_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4152" *)
  wire mux_616_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4151" *)
  wire mux_617_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2858" *)
  wire mux_61_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3309" *)
  wire mux_620_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3308" *)
  wire mux_621_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3307" *)
  wire mux_622_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3314" *)
  wire mux_624_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3317" *)
  wire mux_625_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3313" *)
  wire mux_627_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3319" *)
  wire mux_628_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2863" *)
  wire mux_62_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3318" *)
  wire mux_631_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3312" *)
  wire mux_634_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3327" *)
  wire mux_635_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3330" *)
  wire mux_636_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3326" *)
  wire mux_638_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4157" *)
  wire mux_639_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2862" *)
  wire mux_63_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3325" *)
  wire mux_645_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3333" *)
  wire mux_646_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3336" *)
  wire mux_647_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3332" *)
  wire mux_649_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2867" *)
  wire mux_64_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3331" *)
  wire mux_650_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3324" *)
  wire mux_651_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3338" *)
  wire mux_652_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3337" *)
  wire mux_653_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3341" *)
  wire mux_654_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3344" *)
  wire mux_655_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3347" *)
  wire mux_657_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3350" *)
  wire mux_658_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3353" *)
  wire mux_659_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2866" *)
  wire mux_65_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3355" *)
  wire mux_660_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3358" *)
  wire mux_661_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3365" *)
  wire mux_662_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3363" *)
  wire mux_663_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3370" *)
  wire mux_664_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3373" *)
  wire mux_665_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3369" *)
  wire mux_666_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3361" *)
  wire mux_667_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3376" *)
  wire mux_668_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2861" *)
  wire mux_66_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2549" *)
  wire mux_670_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3377" *)
  wire mux_671_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3378" *)
  wire mux_672_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3383" *)
  wire mux_673_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3381" *)
  wire mux_674_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3388" *)
  wire mux_675_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3390" *)
  wire mux_676_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3387" *)
  wire mux_677_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3379" *)
  wire mux_678_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2875" *)
  wire mux_67_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3397" *)
  wire mux_684_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3395" *)
  wire mux_685_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3402" *)
  wire mux_686_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3404" *)
  wire mux_687_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3401" *)
  wire mux_688_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3393" *)
  wire mux_689_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2877" *)
  wire mux_68_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3411" *)
  wire mux_695_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3409" *)
  wire mux_696_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3416" *)
  wire mux_697_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3418" *)
  wire mux_698_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3415" *)
  wire mux_699_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2874" *)
  wire mux_69_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3407" *)
  wire mux_700_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3421" *)
  wire mux_704_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3423" *)
  wire mux_706_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3422" *)
  wire mux_707_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4135" *)
  wire mux_70_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3427" *)
  wire mux_710_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3425" *)
  wire mux_711_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3429" *)
  wire mux_715_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3430" *)
  wire mux_716_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3428" *)
  wire mux_717_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3433" *)
  wire mux_721_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3431" *)
  wire mux_722_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3434" *)
  wire mux_729_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4137" *)
  wire mux_72_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3436" *)
  wire mux_730_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3438" *)
  wire mux_731_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3435" *)
  wire mux_732_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3439" *)
  wire mux_735_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3441" *)
  wire mux_737_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3442" *)
  wire mux_738_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3440" *)
  wire mux_739_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3444" *)
  wire mux_743_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2551" *)
  wire mux_745_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3448" *)
  wire mux_746_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3447" *)
  wire mux_747_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3446" *)
  wire mux_748_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3445" *)
  wire mux_749_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2881" *)
  wire mux_74_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3452" *)
  wire mux_751_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3449" *)
  wire mux_754_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1946" *)
  wire mux_755_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3456" *)
  wire mux_756_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3455" *)
  wire mux_757_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3454" *)
  wire mux_758_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3450" *)
  wire mux_759_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2880" *)
  wire mux_75_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3460" *)
  wire mux_761_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3463" *)
  wire mux_766_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3462" *)
  wire mux_767_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3458" *)
  wire mux_768_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3466" *)
  wire mux_769_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4139" *)
  wire mux_76_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2552" *)
  wire mux_771_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3471" *)
  wire mux_772_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3470" *)
  wire mux_773_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3469" *)
  wire mux_774_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3468" *)
  wire mux_775_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3482" *)
  wire mux_783_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3485" *)
  wire mux_784_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3488" *)
  wire mux_785_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1937" *)
  wire mux_789_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4141" *)
  wire mux_78_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3506" *)
  wire mux_790_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3505" *)
  wire mux_791_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3504" *)
  wire mux_792_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2585" *)
  wire mux_793_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3509" *)
  wire mux_796_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3508" *)
  wire mux_797_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3510" *)
  wire mux_798_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3511" *)
  wire mux_799_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3522" *)
  wire mux_803_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2590" *)
  wire mux_805_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3523" *)
  wire mux_806_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2884" *)
  wire mux_80_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3526" *)
  wire mux_815_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2883" *)
  wire mux_81_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3529" *)
  wire mux_820_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3528" *)
  wire mux_821_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3527" *)
  wire mux_822_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3524" *)
  wire mux_823_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3533" *)
  wire mux_825_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2879" *)
  wire mux_82_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3536" *)
  wire mux_830_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3535" *)
  wire mux_831_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3531" *)
  wire mux_832_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2560" *)
  wire mux_83_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3543" *)
  wire mux_840_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3546" *)
  wire mux_841_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1938" *)
  wire mux_845_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3562" *)
  wire mux_846_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3561" *)
  wire mux_847_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3560" *)
  wire mux_848_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2887" *)
  wire mux_84_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2670" *)
  wire mux_851_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3565" *)
  wire mux_852_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3564" *)
  wire mux_853_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3566" *)
  wire mux_854_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3567" *)
  wire mux_855_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3572" *)
  wire mux_859_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2888" *)
  wire mux_85_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3574" *)
  wire mux_861_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2886" *)
  wire mux_86_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3577" *)
  wire mux_870_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3580" *)
  wire mux_875_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3579" *)
  wire mux_876_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3578" *)
  wire mux_877_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3575" *)
  wire mux_878_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2893" *)
  wire mux_87_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3584" *)
  wire mux_880_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3587" *)
  wire mux_885_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3586" *)
  wire mux_886_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3582" *)
  wire mux_887_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2892" *)
  wire mux_88_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3594" *)
  wire mux_895_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3597" *)
  wire mux_896_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2889" *)
  wire mux_89_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1939" *)
  wire mux_900_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3613" *)
  wire mux_901_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3612" *)
  wire mux_902_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3611" *)
  wire mux_903_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3615" *)
  wire mux_910_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3616" *)
  wire mux_912_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3622" *)
  wire mux_916_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3625" *)
  wire mux_917_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3626" *)
  wire mux_918_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3624" *)
  wire mux_919_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3627" *)
  wire mux_926_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2899" *)
  wire mux_92_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3637" *)
  wire mux_933_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3636" *)
  wire mux_934_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3635" *)
  wire mux_935_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3631" *)
  wire mux_936_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3644" *)
  wire mux_943_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3643" *)
  wire mux_944_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3639" *)
  wire mux_945_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3675" *)
  wire mux_949_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3646" *)
  wire mux_953_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3655" *)
  wire mux_954_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3658" *)
  wire mux_955_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1940" *)
  wire mux_959_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3673" *)
  wire mux_961_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3672" *)
  wire mux_962_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3676" *)
  wire mux_969_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3677" *)
  wire mux_971_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3683" *)
  wire mux_975_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3686" *)
  wire mux_980_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3684" *)
  wire mux_981_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2539" *)
  wire mux_982_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3690" *)
  wire mux_986_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3691" *)
  wire mux_995_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3697" *)
  wire mux_996_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3695" *)
  wire mux_997_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3725" *)
  wire mux_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1084" *)
  wire mux_tmp_10;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1185" *)
  wire mux_tmp_1101;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1186" *)
  wire mux_tmp_1104;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1202" *)
  wire mux_tmp_1130;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1204" *)
  wire mux_tmp_1136;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1205" *)
  wire mux_tmp_1143;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1207" *)
  wire mux_tmp_1149;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1208" *)
  wire mux_tmp_1156;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1210" *)
  wire mux_tmp_1162;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1211" *)
  wire mux_tmp_1169;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1213" *)
  wire mux_tmp_1175;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2152" *)
  wire mux_tmp_1247;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2154" *)
  wire mux_tmp_1250;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2156" *)
  wire mux_tmp_1253;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2158" *)
  wire mux_tmp_1257;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1102" *)
  wire mux_tmp_128;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1110" *)
  wire mux_tmp_207;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1113" *)
  wire mux_tmp_220;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1126" *)
  wire mux_tmp_265;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1128" *)
  wire mux_tmp_270;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1130" *)
  wire mux_tmp_279;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1131" *)
  wire mux_tmp_281;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1134" *)
  wire mux_tmp_292;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1137" *)
  wire mux_tmp_301;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1087" *)
  wire mux_tmp_35;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1083" *)
  wire mux_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1144" *)
  wire mux_tmp_475;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1149" *)
  wire mux_tmp_595;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1150" *)
  wire mux_tmp_596;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1152" *)
  wire mux_tmp_617;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1153" *)
  wire mux_tmp_618;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1154" *)
  wire mux_tmp_643;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1157" *)
  wire mux_tmp_655;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1095" *)
  wire mux_tmp_70;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1159" *)
  wire mux_tmp_704;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1096" *)
  wire mux_tmp_72;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1098" *)
  wire mux_tmp_76;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1099" *)
  wire mux_tmp_78;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1181" *)
  wire mux_tmp_978;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3620" *)
  wire nand_102_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4206" *)
  wire nand_113_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4208" *)
  wire nand_114_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4213" *)
  wire nand_115_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4215" *)
  wire nand_116_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4220" *)
  wire nand_117_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4222" *)
  wire nand_118_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3315" *)
  wire nand_15_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3328" *)
  wire nand_16_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3334" *)
  wire nand_17_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3389" *)
  wire nand_18_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3403" *)
  wire nand_19_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3417" *)
  wire nand_20_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3826" *)
  wire nand_33_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3032" *)
  wire nand_76_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4143" *)
  wire nand_93_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2530" *)
  wire nand_95_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3681" *)
  wire nand_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1171" *)
  wire nand_tmp_22;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1103" *)
  wire nand_tmp_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4090" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4084" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4086" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4088" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3914" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpAdd_8U_23U_2_is_a_greater_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3916" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpAdd_8U_23U_2_is_a_greater_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3918" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpAdd_8U_23U_2_is_a_greater_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3912" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_FpAdd_8U_23U_2_is_a_greater_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4184" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4186" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4188" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4182" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4098" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4092" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4094" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4096" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 24 25" *)
  wire [25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3516" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1942" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4641" *)
  wire [323:0] nl_NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_inst_chn_lut_out_rsci_d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3278" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3282" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_11_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3266" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3294" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_5_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3270" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_6_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3290" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_7_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3274" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_8_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3286" *)
  (* unused_bits = "0 9" *)
  wire [9:0] nl_acc_9_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4435" *)
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4438" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4429" *)
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4432" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2784" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2786" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4116" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4124" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4452" *)
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4457" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4456" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4441" *)
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a;
  wire [4:0] nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s;
  wire [3:0] nl_lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2794" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2792" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3920" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2873" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3935" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3938" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4423" *)
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4426" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2380" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4417" *)
  wire [23:0] nl_lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4420" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2378" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2788" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2790" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2429" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3929" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl;
  wire [7:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4238" *)
  wire [23:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a;
  wire [8:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4008" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 248" *)
  wire [248:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1064" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4244" *)
  wire [23:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4229" *)
  wire [23:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4232" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4006" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 248" *)
  wire [248:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1066" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4235" *)
  wire [23:0] nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3892" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3889" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4100" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4102" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_lut_lookup_1_FpNormalize_8U_49U_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2871" *)
  (* unused_bits = "8 9" *)
  wire [9:0] nl_lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4606" *)
  wire [48:0] nl_lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2427" *)
  (* unused_bits = "8 9" *)
  wire [9:0] nl_lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4601" *)
  wire [48:0] nl_lut_lookup_1_FpNormalize_8U_49U_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3475" *)
  (* unused_bits = "31" *)
  wire [31:0] nl_lut_lookup_1_IntLog2_32U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4389" *)
  wire [31:0] nl_lut_lookup_1_IntLog2_32U_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4608" *)
  wire [158:0] nl_lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4603" *)
  wire [158:0] nl_lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3880" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_1_else_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3514" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_1_else_1_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2364" *)
  (* unused_bits = "32" *)
  wire [32:0] nl_lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4320" *)
  wire [8:0] nl_lut_lookup_1_else_1_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4076" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_1_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2225" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_1_else_else_else_else_acc_itm_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2362" *)
  (* unused_bits = "32" *)
  wire [32:0] nl_lut_lookup_1_else_else_else_else_le_data_f_acc_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4313" *)
  wire [34:0] nl_lut_lookup_1_else_else_else_else_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4316" *)
  wire [8:0] nl_lut_lookup_1_else_else_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3846" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_1_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4000" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_1_else_if_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3844" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_lut_lookup_1_if_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3860" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_1_if_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3493" *)
  (* unused_bits = "7" *)
  wire [7:0] nl_lut_lookup_1_if_else_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4307" *)
  wire [30:0] nl_lut_lookup_1_if_else_else_else_else_else_rshift_rg_a;
  wire [6:0] nl_lut_lookup_1_if_else_else_else_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3495" *)
  (* unused_bits = "4" *)
  wire [4:0] nl_lut_lookup_1_if_else_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4301" *)
  wire [30:0] nl_lut_lookup_1_if_else_else_else_else_if_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4304" *)
  wire [5:0] nl_lut_lookup_1_if_else_else_else_else_if_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3862" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_1_if_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3992" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 10" *)
  wire [10:0] nl_lut_lookup_1_if_if_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4068" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_1_if_if_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4403" *)
  wire [48:0] nl_lut_lookup_1_leading_sign_49_0_2_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4401" *)
  wire [48:0] nl_lut_lookup_1_leading_sign_49_0_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4481" *)
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4484" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4475" *)
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4478" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2796" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2798" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4118" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4126" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4498" *)
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4503" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4502" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4487" *)
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4492" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4491" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2806" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2804" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3922" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2929" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3951" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3954" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4469" *)
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4472" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2384" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4463" *)
  wire [23:0] nl_lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4466" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2382" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2800" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2802" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2422" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3945" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl;
  wire [7:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4256" *)
  wire [23:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a;
  wire [8:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4019" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 248" *)
  wire [248:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1060" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4262" *)
  wire [23:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4247" *)
  wire [23:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4250" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4017" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 248" *)
  wire [248:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1062" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4253" *)
  wire [23:0] nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3898" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3895" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4104" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4106" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_lut_lookup_2_FpNormalize_8U_49U_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2927" *)
  (* unused_bits = "8 9" *)
  wire [9:0] nl_lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4616" *)
  wire [48:0] nl_lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2420" *)
  (* unused_bits = "8 9" *)
  wire [9:0] nl_lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4611" *)
  wire [48:0] nl_lut_lookup_2_FpNormalize_8U_49U_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3540" *)
  (* unused_bits = "31" *)
  wire [31:0] nl_lut_lookup_2_IntLog2_32U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4392" *)
  wire [31:0] nl_lut_lookup_2_IntLog2_32U_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4618" *)
  wire [158:0] nl_lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4613" *)
  wire [158:0] nl_lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3882" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_2_else_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4342" *)
  wire [8:0] nl_lut_lookup_2_else_1_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4080" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_2_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4335" *)
  wire [34:0] nl_lut_lookup_2_else_else_else_else_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4338" *)
  wire [8:0] nl_lut_lookup_2_else_else_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3850" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_2_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4011" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_2_else_if_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3848" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_lut_lookup_2_if_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3864" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_2_if_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3549" *)
  (* unused_bits = "7" *)
  wire [7:0] nl_lut_lookup_2_if_else_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4329" *)
  wire [30:0] nl_lut_lookup_2_if_else_else_else_else_else_rshift_rg_a;
  wire [6:0] nl_lut_lookup_2_if_else_else_else_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3551" *)
  (* unused_bits = "4" *)
  wire [4:0] nl_lut_lookup_2_if_else_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4323" *)
  wire [30:0] nl_lut_lookup_2_if_else_else_else_else_if_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4326" *)
  wire [5:0] nl_lut_lookup_2_if_else_else_else_else_if_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3866" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_2_if_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3994" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 10" *)
  wire [10:0] nl_lut_lookup_2_if_if_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4070" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_2_if_if_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4407" *)
  wire [48:0] nl_lut_lookup_2_leading_sign_49_0_2_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4405" *)
  wire [48:0] nl_lut_lookup_2_leading_sign_49_0_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4527" *)
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4530" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4521" *)
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4524" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2808" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2810" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4120" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4128" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4544" *)
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4549" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4548" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4533" *)
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4538" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4537" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2818" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2816" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3924" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2979" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3967" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3970" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4515" *)
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4518" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2388" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4509" *)
  wire [23:0] nl_lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4512" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2386" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2812" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2814" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2415" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3961" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl;
  wire [7:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4274" *)
  wire [23:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a;
  wire [8:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4030" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 248" *)
  wire [248:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1056" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4280" *)
  wire [23:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4265" *)
  wire [23:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4268" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4028" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 248" *)
  wire [248:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1058" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4271" *)
  wire [23:0] nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3904" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3901" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4108" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4110" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_lut_lookup_3_FpNormalize_8U_49U_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2977" *)
  (* unused_bits = "8 9" *)
  wire [9:0] nl_lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4626" *)
  wire [48:0] nl_lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2413" *)
  (* unused_bits = "8 9" *)
  wire [9:0] nl_lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4621" *)
  wire [48:0] nl_lut_lookup_3_FpNormalize_8U_49U_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3591" *)
  (* unused_bits = "31" *)
  wire [31:0] nl_lut_lookup_3_IntLog2_32U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4395" *)
  wire [31:0] nl_lut_lookup_3_IntLog2_32U_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4628" *)
  wire [158:0] nl_lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4623" *)
  wire [158:0] nl_lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3884" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_3_else_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4364" *)
  wire [8:0] nl_lut_lookup_3_else_1_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4078" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_3_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4357" *)
  wire [34:0] nl_lut_lookup_3_else_else_else_else_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4360" *)
  wire [8:0] nl_lut_lookup_3_else_else_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3854" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_3_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4022" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_3_else_if_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3852" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_lut_lookup_3_if_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3868" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_3_if_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3600" *)
  (* unused_bits = "7" *)
  wire [7:0] nl_lut_lookup_3_if_else_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4351" *)
  wire [30:0] nl_lut_lookup_3_if_else_else_else_else_else_rshift_rg_a;
  wire [6:0] nl_lut_lookup_3_if_else_else_else_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3602" *)
  (* unused_bits = "4" *)
  wire [4:0] nl_lut_lookup_3_if_else_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4345" *)
  wire [30:0] nl_lut_lookup_3_if_else_else_else_else_if_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4348" *)
  wire [5:0] nl_lut_lookup_3_if_else_else_else_else_if_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3870" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_3_if_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3996" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 10" *)
  wire [10:0] nl_lut_lookup_3_if_if_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4072" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_3_if_if_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4411" *)
  wire [48:0] nl_lut_lookup_3_leading_sign_49_0_2_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4409" *)
  wire [48:0] nl_lut_lookup_3_leading_sign_49_0_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4573" *)
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4576" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4567" *)
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4570" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2820" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2822" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4122" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4130" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4590" *)
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4595" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4594" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4579" *)
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4584" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4583" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2830" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2828" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3926" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3029" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3983" *)
  (* unused_bits = "0 1 2 3 4 5 6 8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3986" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4561" *)
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4564" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2392" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4555" *)
  wire [23:0] nl_lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4558" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2390" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2824" *)
  (* unused_bits = "50 51" *)
  wire [51:0] nl_lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2826" *)
  (* unused_bits = "50" *)
  wire [50:0] nl_lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2408" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3977" *)
  (* unused_bits = "8" *)
  wire [8:0] nl_lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl;
  wire [7:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4292" *)
  wire [23:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a;
  wire [8:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4041" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 248" *)
  wire [248:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1052" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4298" *)
  wire [23:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4283" *)
  wire [23:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a;
  wire [7:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4039" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 248" *)
  wire [248:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1054" *)
  (* unused_bits = "10" *)
  wire [10:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4289" *)
  wire [23:0] nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3910" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3907" *)
  (* unused_bits = "23" *)
  wire [23:0] nl_lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4112" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4114" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 9 10" *)
  wire [10:0] nl_lut_lookup_4_FpNormalize_8U_49U_2_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3027" *)
  (* unused_bits = "8 9" *)
  wire [9:0] nl_lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4636" *)
  wire [48:0] nl_lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2406" *)
  (* unused_bits = "8 9" *)
  wire [9:0] nl_lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4631" *)
  wire [48:0] nl_lut_lookup_4_FpNormalize_8U_49U_else_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3652" *)
  (* unused_bits = "31" *)
  wire [31:0] nl_lut_lookup_4_IntLog2_32U_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4398" *)
  wire [31:0] nl_lut_lookup_4_IntLog2_32U_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4638" *)
  wire [158:0] nl_lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4633" *)
  wire [158:0] nl_lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3886" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_4_else_1_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4386" *)
  wire [8:0] nl_lut_lookup_4_else_1_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4082" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_4_else_else_acc_1_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4379" *)
  wire [34:0] nl_lut_lookup_4_else_else_else_else_rshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4382" *)
  wire [8:0] nl_lut_lookup_4_else_else_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3858" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_4_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4033" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_4_else_if_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3856" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 11" *)
  wire [11:0] nl_lut_lookup_4_if_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3872" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 33" *)
  wire [33:0] nl_lut_lookup_4_if_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3661" *)
  (* unused_bits = "7" *)
  wire [7:0] nl_lut_lookup_4_if_else_else_else_else_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4373" *)
  wire [30:0] nl_lut_lookup_4_if_else_else_else_else_else_rshift_rg_a;
  wire [6:0] nl_lut_lookup_4_if_else_else_else_else_else_rshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3663" *)
  (* unused_bits = "4" *)
  wire [4:0] nl_lut_lookup_4_if_else_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4367" *)
  wire [30:0] nl_lut_lookup_4_if_else_else_else_else_if_lshift_rg_a;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4370" *)
  wire [5:0] nl_lut_lookup_4_if_else_else_else_else_if_lshift_rg_s;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3874" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_4_if_else_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3998" *)
  (* unused_bits = "0 1 2 3 4 5 6 7 8 10" *)
  wire [10:0] nl_lut_lookup_4_if_if_else_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4074" *)
  (* unused_bits = "0 1 2 4" *)
  wire [4:0] nl_lut_lookup_4_if_if_else_else_if_acc_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4415" *)
  wire [48:0] nl_lut_lookup_4_leading_sign_49_0_2_rg_mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4413" *)
  wire [48:0] nl_lut_lookup_4_leading_sign_49_0_rg_mantissa;
  wire [31:0] nl_lut_lookup_else_1_lo_index_u_1_sva_3;
  wire [31:0] nl_lut_lookup_else_1_lo_index_u_2_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1536" *)
  (* unused_bits = "32" *)
  wire [32:0] nl_lut_lookup_else_1_lo_index_u_3_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1566" *)
  (* unused_bits = "32" *)
  wire [32:0] nl_lut_lookup_else_1_lo_index_u_sva_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1952" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_if_else_else_else_le_index_s_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1954" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_if_else_else_else_le_index_s_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1956" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_if_else_else_else_le_index_s_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1958" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_if_else_else_else_le_index_s_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2211" *)
  (* unused_bits = "32" *)
  wire [32:0] nl_lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2213" *)
  (* unused_bits = "32" *)
  wire [32:0] nl_lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2215" *)
  (* unused_bits = "32" *)
  wire [32:0] nl_lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2217" *)
  (* unused_bits = "32" *)
  wire [32:0] nl_lut_lookup_if_else_else_le_data_sub_sva_mx0w0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1825" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_if_if_else_else_le_index_s_1_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1823" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_if_if_else_else_le_index_s_2_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1821" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_if_if_else_else_le_index_s_3_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1819" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_lut_lookup_if_if_else_else_le_index_s_sva;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2162" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_z_out_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2164" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_z_out_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2166" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_z_out_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2168" *)
  (* unused_bits = "9" *)
  wire [9:0] nl_z_out_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1849" *)
  wire nor_13_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2527" *)
  wire nor_190_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2542" *)
  wire nor_193_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2448" *)
  wire nor_27_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1850" *)
  wire nor_31_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2453" *)
  wire nor_38_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3668" *)
  wire nor_412_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3669" *)
  wire nor_413_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3665" *)
  wire nor_414_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3666" *)
  wire nor_415_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3607" *)
  wire nor_418_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3608" *)
  wire nor_419_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3604" *)
  wire nor_420_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3605" *)
  wire nor_421_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3556" *)
  wire nor_424_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3557" *)
  wire nor_425_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3553" *)
  wire nor_426_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3554" *)
  wire nor_427_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1851" *)
  wire nor_42_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3500" *)
  wire nor_430_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3501" *)
  wire nor_431_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3497" *)
  wire nor_432_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3498" *)
  wire nor_433_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3490" *)
  wire nor_434_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3491" *)
  wire nor_435_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4179" *)
  wire nor_438_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4176" *)
  wire nor_440_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4173" *)
  wire nor_442_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4170" *)
  wire nor_444_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3838" *)
  wire nor_448_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3839" *)
  wire nor_449_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3835" *)
  wire nor_450_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3831" *)
  wire nor_451_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3815" *)
  wire nor_453_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3818" *)
  wire nor_454_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3804" *)
  wire nor_455_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3793" *)
  wire nor_459_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3781" *)
  wire nor_463_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3784" *)
  wire nor_464_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3775" *)
  wire nor_465_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3776" *)
  wire nor_466_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3772" *)
  wire nor_467_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3773" *)
  wire nor_468_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1881" *)
  wire nor_469_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3769" *)
  wire nor_470_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3770" *)
  wire nor_471_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3766" *)
  wire nor_472_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3767" *)
  wire nor_473_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3761" *)
  wire nor_475_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3763" *)
  wire nor_476_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3764" *)
  wire nor_477_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3758" *)
  wire nor_478_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3759" *)
  wire nor_479_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3755" *)
  wire nor_480_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3756" *)
  wire nor_481_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1882" *)
  wire nor_482_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3752" *)
  wire nor_483_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3753" *)
  wire nor_484_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3749" *)
  wire nor_485_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3750" *)
  wire nor_486_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3746" *)
  wire nor_487_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3747" *)
  wire nor_488_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3743" *)
  wire nor_489_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3744" *)
  wire nor_490_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3740" *)
  wire nor_491_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3741" *)
  wire nor_492_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3737" *)
  wire nor_493_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3738" *)
  wire nor_494_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3732" *)
  wire nor_495_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3734" *)
  wire nor_496_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3735" *)
  wire nor_497_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3718" *)
  wire nor_500_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3720" *)
  wire nor_501_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3721" *)
  wire nor_503_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3708" *)
  wire nor_506_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3710" *)
  wire nor_507_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3711" *)
  wire nor_509_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2456" *)
  wire nor_50_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3696" *)
  wire nor_512_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3698" *)
  wire nor_513_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3699" *)
  wire nor_515_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3685" *)
  wire nor_518_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3687" *)
  wire nor_519_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3688" *)
  wire nor_521_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1895" *)
  wire nor_526_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3656" *)
  wire nor_528_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3657" *)
  wire nor_529_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3634" *)
  wire nor_540_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3630" *)
  wire nor_544_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3614" *)
  wire nor_549_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1852" *)
  wire nor_54_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3595" *)
  wire nor_551_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3596" *)
  wire nor_552_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1949" *)
  wire nor_564_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3563" *)
  wire nor_573_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3544" *)
  wire nor_575_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3545" *)
  wire nor_576_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1948" *)
  wire nor_588_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3507" *)
  wire nor_595_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3483" *)
  wire nor_597_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3484" *)
  wire nor_598_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2442" *)
  wire nor_5_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3467" *)
  wire nor_606_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3472" *)
  wire nor_609_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1894" *)
  wire nor_610_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1870" *)
  wire nor_612_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3453" *)
  wire nor_616_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3437" *)
  wire nor_619_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4160" *)
  wire nor_622_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3412" *)
  wire nor_623_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3419" *)
  wire nor_626_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3398" *)
  wire nor_628_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3405" *)
  wire nor_631_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3384" *)
  wire nor_633_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2567" *)
  wire nor_634_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3391" *)
  wire nor_636_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3366" *)
  wire nor_638_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3374" *)
  wire nor_640_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4159" *)
  wire nor_641_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3339" *)
  wire nor_642_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4155" *)
  wire nor_647_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3245" *)
  wire nor_657_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3231" *)
  wire nor_658_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3232" *)
  wire nor_659_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3228" *)
  wire nor_660_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3229" *)
  wire nor_661_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3223" *)
  wire nor_662_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3224" *)
  wire nor_663_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3220" *)
  wire nor_664_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3221" *)
  wire nor_665_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3205" *)
  wire nor_666_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3206" *)
  wire nor_667_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3199" *)
  wire nor_668_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3200" *)
  wire nor_669_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3194" *)
  wire nor_670_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3195" *)
  wire nor_671_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3191" *)
  wire nor_672_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3192" *)
  wire nor_673_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3182" *)
  wire nor_674_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3183" *)
  wire nor_675_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3179" *)
  wire nor_676_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3180" *)
  wire nor_677_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3170" *)
  wire nor_678_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3172" *)
  wire nor_679_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3173" *)
  wire nor_680_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3165" *)
  wire nor_681_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3167" *)
  wire nor_682_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3168" *)
  wire nor_683_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3162" *)
  wire nor_684_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3163" *)
  wire nor_685_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3159" *)
  wire nor_686_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3160" *)
  wire nor_687_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3150" *)
  wire nor_689_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2668" *)
  wire nor_690_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3148" *)
  wire nor_691_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3145" *)
  wire nor_692_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3146" *)
  wire nor_693_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3137" *)
  wire nor_694_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3138" *)
  wire nor_695_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3132" *)
  wire nor_696_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3133" *)
  wire nor_697_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3129" *)
  wire nor_698_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3130" *)
  wire nor_699_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3120" *)
  wire nor_700_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3113" *)
  wire nor_701_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3114" *)
  wire nor_702_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3110" *)
  wire nor_705_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3111" *)
  wire nor_706_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3093" *)
  wire nor_707_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3094" *)
  wire nor_708_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3090" *)
  wire nor_711_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3091" *)
  wire nor_712_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3076" *)
  wire nor_713_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3079" *)
  wire nor_714_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3072" *)
  wire nor_715_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3073" *)
  wire nor_716_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3069" *)
  wire nor_719_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3070" *)
  wire nor_720_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3057" *)
  wire nor_721_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3050" *)
  wire nor_722_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3051" *)
  wire nor_723_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3047" *)
  wire nor_724_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3048" *)
  wire nor_725_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3044" *)
  wire nor_726_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3045" *)
  wire nor_727_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3020" *)
  wire nor_729_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3024" *)
  wire nor_730_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3015" *)
  wire nor_732_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3016" *)
  wire nor_733_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2999" *)
  wire nor_737_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3000" *)
  wire nor_738_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2970" *)
  wire nor_742_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2974" *)
  wire nor_743_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2965" *)
  wire nor_745_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2966" *)
  wire nor_746_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2949" *)
  wire nor_749_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2950" *)
  wire nor_750_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2920" *)
  wire nor_757_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2924" *)
  wire nor_758_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2915" *)
  wire nor_760_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2916" *)
  wire nor_761_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2900" *)
  wire nor_764_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2901" *)
  wire nor_765_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2864" *)
  wire nor_769_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2868" *)
  wire nor_770_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2859" *)
  wire nor_772_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2860" *)
  wire nor_773_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2842" *)
  wire nor_775_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2843" *)
  wire nor_776_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4133" *)
  wire nor_779_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2782" *)
  wire nor_783_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2484" *)
  wire nor_792_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2499" *)
  wire nor_813_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4201" *)
  wire nor_814_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4197" *)
  wire nor_817_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4196" *)
  wire nor_820_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4195" *)
  wire nor_823_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3680" *)
  wire nor_825_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3619" *)
  wire nor_827_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3520" *)
  wire nor_830_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3479" *)
  wire nor_831_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2493" *)
  wire nor_832_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3481" *)
  wire nor_833_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2908" *)
  wire nor_852_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2508" *)
  wire nor_855_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2523" *)
  wire nor_865_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2438" *)
  wire nor_874_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3117" *)
  wire nor_879_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3097" *)
  wire nor_880_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3054" *)
  wire nor_881_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4227" *)
  wire nor_882_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1143" *)
  wire nor_tmp_112;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1092" *)
  wire nor_tmp_12;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1093" *)
  wire nor_tmp_14;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1165" *)
  wire nor_tmp_238;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1170" *)
  wire nor_tmp_260;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1174" *)
  wire nor_tmp_281;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1100" *)
  wire nor_tmp_32;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1101" *)
  wire nor_tmp_34;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1105" *)
  wire nor_tmp_44;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1106" *)
  wire nor_tmp_46;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1108" *)
  wire nor_tmp_55;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1109" *)
  wire nor_tmp_57;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1112" *)
  wire not_tmp_209;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1116" *)
  wire not_tmp_222;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1118" *)
  wire not_tmp_235;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1123" *)
  wire not_tmp_248;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1133" *)
  wire not_tmp_276;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1142" *)
  wire not_tmp_334;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1145" *)
  wire not_tmp_394;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1146" *)
  wire not_tmp_412;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1147" *)
  wire not_tmp_418;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1148" *)
  wire not_tmp_422;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1085" *)
  wire not_tmp_47;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1183" *)
  wire not_tmp_800;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:938" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:939" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3512" *)
  wire or_1045_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3530" *)
  wire or_1072_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3568" *)
  wire or_1113_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3581" *)
  wire or_1142_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2876" *)
  wire or_114_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3617" *)
  wire or_1183_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2878" *)
  wire or_118_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1900" *)
  wire or_1202_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2882" *)
  wire or_120_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3638" *)
  wire or_1213_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4138" *)
  wire or_121_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4136" *)
  wire or_122_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3678" *)
  wire or_1252_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2885" *)
  wire or_125_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4142" *)
  wire or_126_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4140" *)
  wire or_127_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3788" *)
  wire or_1431_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3799" *)
  wire or_1440_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3810" *)
  wire or_1450_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3822" *)
  wire or_1458_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3828" *)
  wire or_1460_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1905" *)
  wire or_1495_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4162" *)
  wire or_1583_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4164" *)
  wire or_1594_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4166" *)
  wire or_1606_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4168" *)
  wire or_1618_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2529" *)
  wire or_1688_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1891" *)
  wire or_1689_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2538" *)
  wire or_1691_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3322" *)
  wire or_1696_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3827" *)
  wire or_1830_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2933" *)
  wire or_184_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2584" *)
  wire or_1851_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1864" *)
  wire or_1853_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1868" *)
  wire or_1857_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4150" *)
  wire or_1860_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4145" *)
  wire or_186_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4144" *)
  wire or_191_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2839" *)
  wire or_1931_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2520" *)
  wire or_1936_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2850" *)
  wire or_1941_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2897" *)
  wire or_1948_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2946" *)
  wire or_1964_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4190" *)
  wire or_1972_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4191" *)
  wire or_1973_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2956" *)
  wire or_1976_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2996" *)
  wire or_1983_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4193" *)
  wire or_1991_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4194" *)
  wire or_1992_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3006" *)
  wire or_1995_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3521" *)
  wire or_2007_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3518" *)
  wire or_2009_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3621" *)
  wire or_2025_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3682" *)
  wire or_2035_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4200" *)
  wire or_2055_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4199" *)
  wire or_2056_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2994" *)
  wire or_2078_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2944" *)
  wire or_2079_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2895" *)
  wire or_2080_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2837" *)
  wire or_2081_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3649" *)
  wire or_2087_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4207" *)
  wire or_2088_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4214" *)
  wire or_2089_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4221" *)
  wire or_2090_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2982" *)
  wire or_247_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2984" *)
  wire or_251_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1866" *)
  wire or_26_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4146" *)
  wire or_302_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3034" *)
  wire or_306_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3040" *)
  wire or_311_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2547" *)
  wire or_312_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3042" *)
  wire or_315_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3059" *)
  wire or_332_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3065" *)
  wire or_341_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3067" *)
  wire or_346_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2669" *)
  wire or_365_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3086" *)
  wire or_374_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3106" *)
  wire or_406_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2891" *)
  wire or_40_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3108" *)
  wire or_411_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3135" *)
  wire or_445_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3152" *)
  wire or_475_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2498" *)
  wire or_48_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2565" *)
  wire or_492_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4131" *)
  wire or_4_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3186" *)
  wire or_528_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3197" *)
  wire or_545_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3208" *)
  wire or_566_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3210" *)
  wire or_569_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3212" *)
  wire or_575_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3226" *)
  wire or_596_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3234" *)
  wire or_617_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3236" *)
  wire or_620_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3238" *)
  wire or_625_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1873" *)
  wire or_66_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3302" *)
  wire or_827_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3306" *)
  wire or_829_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4156" *)
  wire or_832_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3311" *)
  wire or_839_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4154" *)
  wire or_841_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2526" *)
  wire or_849_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3320" *)
  wire or_850_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4158" *)
  wire or_856_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3364" *)
  wire or_879_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3367" *)
  wire or_880_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3371" *)
  wire or_885_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3372" *)
  wire or_887_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3375" *)
  wire or_888_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3382" *)
  wire or_899_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3385" *)
  wire or_900_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3392" *)
  wire or_907_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3396" *)
  wire or_915_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3399" *)
  wire or_916_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3406" *)
  wire or_923_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3410" *)
  wire or_931_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3413" *)
  wire or_932_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3420" *)
  wire or_939_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1880" *)
  wire or_969_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1869" *)
  wire or_978_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:3457" *)
  wire or_990_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2435" *)
  wire or_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1198" *)
  wire or_dcpl_51;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1201" *)
  wire or_dcpl_57;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1091" *)
  wire or_tmp_101;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1167" *)
  wire or_tmp_1043;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1175" *)
  wire or_tmp_1181;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1094" *)
  wire or_tmp_124;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1179" *)
  wire or_tmp_1250;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1097" *)
  wire or_tmp_129;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1182" *)
  wire or_tmp_1360;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1184" *)
  wire or_tmp_1450;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1195" *)
  wire or_tmp_1490;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1203" *)
  wire or_tmp_1513;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1206" *)
  wire or_tmp_1523;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1209" *)
  wire or_tmp_1534;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1212" *)
  wire or_tmp_1545;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1232" *)
  wire or_tmp_1628;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1982" *)
  wire or_tmp_1663;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1984" *)
  wire or_tmp_1671;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1989" *)
  wire or_tmp_1674;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1990" *)
  wire or_tmp_1678;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1994" *)
  wire or_tmp_1684;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1995" *)
  wire or_tmp_1692;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1999" *)
  wire or_tmp_1697;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2000" *)
  wire or_tmp_1705;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2001" *)
  wire or_tmp_1707;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2043" *)
  wire or_tmp_1716;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2046" *)
  wire or_tmp_1720;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1111" *)
  wire or_tmp_314;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1114" *)
  wire or_tmp_331;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1117" *)
  wire or_tmp_363;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1119" *)
  wire or_tmp_378;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1120" *)
  wire or_tmp_380;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1121" *)
  wire or_tmp_395;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1122" *)
  wire or_tmp_397;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1124" *)
  wire or_tmp_427;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1125" *)
  wire or_tmp_428;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1086" *)
  wire or_tmp_44;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1127" *)
  wire or_tmp_447;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1129" *)
  wire or_tmp_456;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1132" *)
  wire or_tmp_478;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1135" *)
  wire or_tmp_505;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1136" *)
  wire or_tmp_522;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1138" *)
  wire or_tmp_547;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1139" *)
  wire or_tmp_573;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1140" *)
  wire or_tmp_598;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1081" *)
  wire or_tmp_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1141" *)
  wire or_tmp_623;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1088" *)
  wire or_tmp_63;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1082" *)
  wire or_tmp_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1151" *)
  wire or_tmp_843;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1161" *)
  wire or_tmp_976;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1162" *)
  wire or_tmp_980;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1163" *)
  wire or_tmp_993;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2067" *)
  reg [5:0] reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2066" *)
  reg [1:0] reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2071" *)
  reg [5:0] reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2070" *)
  reg [1:0] reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2075" *)
  reg [5:0] reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2074" *)
  reg [1:0] reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2079" *)
  reg [5:0] reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2078" *)
  reg [1:0] reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2054" *)
  reg [5:0] reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2053" *)
  reg [1:0] reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2057" *)
  reg [5:0] reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2056" *)
  reg [1:0] reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2060" *)
  reg [5:0] reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2059" *)
  reg [1:0] reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2063" *)
  reg [5:0] reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2062" *)
  reg [1:0] reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2115" *)
  reg [22:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2114" *)
  reg [7:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1920" *)
  reg [22:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1919" *)
  reg [7:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1932" *)
  reg [22:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1926" *)
  reg [22:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1925" *)
  reg [7:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1931" *)
  reg [7:0] reg_IntLog2_32U_ac_int_cctor_1_30_0_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2543" *)
  reg reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2558" *)
  reg reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2505" *)
  reg reg_cfg_lut_le_function_1_sva_st_19_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2522" *)
  reg reg_cfg_lut_le_function_1_sva_st_20_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2504" *)
  reg [1:0] reg_cfg_precision_1_sva_st_12_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2521" *)
  reg [1:0] reg_cfg_precision_1_sva_st_13_cse_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1865" *)
  reg reg_chn_lut_out_rsci_ld_core_psct_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2510" *)
  reg reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2511" *)
  reg reg_lut_lookup_1_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2445" *)
  reg reg_lut_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2118" *)
  reg [7:0] reg_lut_lookup_1_else_1_else_else_acc_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2117" *)
  reg reg_lut_lookup_1_else_1_else_else_acc_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1916" *)
  reg reg_lut_lookup_1_else_else_else_else_acc_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1917" *)
  reg [2:0] reg_lut_lookup_1_else_else_else_else_acc_2_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1918" *)
  reg [3:0] reg_lut_lookup_1_else_else_else_else_acc_3_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1915" *)
  reg reg_lut_lookup_1_else_else_else_else_acc_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2065" *)
  reg [1:0] reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2064" *)
  reg reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2512" *)
  reg reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2475" *)
  reg reg_lut_lookup_2_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2450" *)
  reg reg_lut_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2121" *)
  reg [7:0] reg_lut_lookup_2_else_1_else_else_acc_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2120" *)
  reg reg_lut_lookup_2_else_1_else_else_acc_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1922" *)
  reg reg_lut_lookup_2_else_else_else_else_acc_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1923" *)
  reg [2:0] reg_lut_lookup_2_else_else_else_else_acc_2_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1924" *)
  reg [3:0] reg_lut_lookup_2_else_else_else_else_acc_3_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1921" *)
  reg reg_lut_lookup_2_else_else_else_else_acc_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2069" *)
  reg [1:0] reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2068" *)
  reg reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2513" *)
  reg reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2514" *)
  reg reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2454" *)
  reg reg_lut_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2124" *)
  reg [7:0] reg_lut_lookup_3_else_1_else_else_acc_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2123" *)
  reg reg_lut_lookup_3_else_1_else_else_acc_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1928" *)
  reg reg_lut_lookup_3_else_else_else_else_acc_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1929" *)
  reg [2:0] reg_lut_lookup_3_else_else_else_else_acc_2_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1930" *)
  reg [3:0] reg_lut_lookup_3_else_else_else_else_acc_3_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1927" *)
  reg reg_lut_lookup_3_else_else_else_else_acc_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2073" *)
  reg [1:0] reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2072" *)
  reg reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2515" *)
  reg reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2516" *)
  reg reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2457" *)
  reg reg_lut_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2127" *)
  reg [7:0] reg_lut_lookup_4_else_1_else_else_acc_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2126" *)
  reg reg_lut_lookup_4_else_1_else_else_acc_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1934" *)
  reg reg_lut_lookup_4_else_else_else_else_acc_1_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1935" *)
  reg [2:0] reg_lut_lookup_4_else_else_else_else_acc_2_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1936" *)
  reg [3:0] reg_lut_lookup_4_else_else_else_else_acc_3_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:1933" *)
  reg reg_lut_lookup_4_else_else_else_else_acc_reg;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2077" *)
  reg [1:0] reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2076" *)
  reg reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2509" *)
  reg reg_lut_lookup_if_unequal_cse;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2153" *)
  wire z_out;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2155" *)
  wire z_out_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2157" *)
  wire z_out_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2160" *)
  wire z_out_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2161" *)
  wire [8:0] z_out_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2163" *)
  wire [8:0] z_out_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2165" *)
  wire [8:0] z_out_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:2167" *)
  wire [8:0] z_out_7;
  assign acc_6_nl = { FpAdd_8U_23U_2_a_right_shift_qelse_mux_10_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11926" *) { FpAdd_8U_23U_2_a_right_shift_qelse_mux_11_nl, 1'b1 };
  assign acc_8_nl = { FpAdd_8U_23U_a_right_shift_qelse_mux_12_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11933" *) { FpAdd_8U_23U_a_right_shift_qelse_mux_13_nl, 1'b1 };
  assign acc_11_nl = { FpAdd_8U_23U_a_right_shift_qelse_mux_14_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11940" *) { FpAdd_8U_23U_a_right_shift_qelse_mux_15_nl, 1'b1 };
  assign acc_7_nl = { FpAdd_8U_23U_a_right_shift_qelse_mux_10_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11947" *) { FpAdd_8U_23U_a_right_shift_qelse_mux_11_nl, 1'b1 };
  assign _00870_ = { 1'b1, _02156_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11950" *) FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0;
  assign lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl = _00870_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11950" *) 1'b1;
  assign lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl = FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11953" *) FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0;
  assign _00871_ = { 1'b1, _02157_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11956" *) FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0;
  assign lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl = _00871_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11956" *) 1'b1;
  assign lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl = FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11959" *) FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0;
  assign lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl = FpAdd_8U_23U_2_addend_larger_qr_1_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11962" *) FpAdd_8U_23U_2_addend_smaller_qr_1_lpi_1_dfm_mx0;
  assign _00872_ = { 1'b1, _02158_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11965" *) FpAdd_8U_23U_2_addend_larger_qr_1_lpi_1_dfm_mx0;
  assign lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl = _00872_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11965" *) 1'b1;
  assign _00873_ = { 1'b1, _02159_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11968" *) FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0;
  assign lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl = _00873_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11968" *) 1'b1;
  assign lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl = FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11971" *) FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0;
  assign _00874_ = { 1'b1, _02160_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11974" *) FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0;
  assign lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl = _00874_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11974" *) 1'b1;
  assign lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl = FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11977" *) FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0;
  assign lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl = FpAdd_8U_23U_2_addend_larger_qr_2_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11980" *) FpAdd_8U_23U_2_addend_smaller_qr_2_lpi_1_dfm_mx0;
  assign _00875_ = { 1'b1, _02161_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11983" *) FpAdd_8U_23U_2_addend_larger_qr_2_lpi_1_dfm_mx0;
  assign lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl = _00875_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11983" *) 1'b1;
  assign _00876_ = { 1'b1, _02162_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11986" *) FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0;
  assign lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl = _00876_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11986" *) 1'b1;
  assign lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl = FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11989" *) FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0;
  assign _00877_ = { 1'b1, _02163_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11992" *) FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0;
  assign lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl = _00877_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11992" *) 1'b1;
  assign lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl = FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11995" *) FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0;
  assign lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl = FpAdd_8U_23U_2_addend_larger_qr_3_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11998" *) FpAdd_8U_23U_2_addend_smaller_qr_3_lpi_1_dfm_mx0;
  assign _00878_ = { 1'b1, _02164_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12001" *) FpAdd_8U_23U_2_addend_larger_qr_3_lpi_1_dfm_mx0;
  assign lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl = _00878_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12001" *) 1'b1;
  assign _00879_ = { 1'b1, _02165_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12004" *) FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0;
  assign lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl = _00879_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12004" *) 1'b1;
  assign lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl = FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12007" *) FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0;
  assign _00880_ = { 1'b1, _02166_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12010" *) FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0;
  assign lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl = _00880_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12010" *) 1'b1;
  assign lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl = FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12013" *) FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0;
  assign lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl = FpAdd_8U_23U_2_addend_larger_qr_lpi_1_dfm_mx0 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12016" *) FpAdd_8U_23U_2_addend_smaller_qr_lpi_1_dfm_mx0;
  assign _00881_ = { 1'b1, _02167_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12019" *) FpAdd_8U_23U_2_addend_larger_qr_lpi_1_dfm_mx0;
  assign lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl = _00881_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12019" *) 1'b1;
  assign _00882_ = FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12067" *) { 2'b11, _02172_ };
  assign lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl = _00882_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12067" *) 1'b1;
  assign lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl = FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12072" *) 1'b1;
  assign _00883_ = FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12135" *) { 2'b11, _02177_ };
  assign lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl = _00883_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12135" *) 1'b1;
  assign lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl = FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12140" *) 1'b1;
  assign _00884_ = FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12197" *) { 2'b11, _02182_ };
  assign lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl = _00884_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12197" *) 1'b1;
  assign lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl = FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12202" *) 1'b1;
  assign _00885_ = FpAdd_8U_23U_2_qr_lpi_1_dfm_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12263" *) { 2'b11, _02186_ };
  assign lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl = _00885_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12263" *) 1'b1;
  assign lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl = FpAdd_8U_23U_2_qr_lpi_1_dfm_5 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12268" *) 1'b1;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_2_tmp + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12297" *) 8'b10000001;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_5_tmp + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12318" *) 8'b10000001;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_8_tmp + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12337" *) 8'b10000001;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_11_tmp + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12358" *) 8'b10000001;
  assign acc_4_nl = { FpAdd_8U_23U_a_right_shift_qelse_mux_8_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12589" *) { FpAdd_8U_23U_a_right_shift_qelse_mux_9_nl, 1'b1 };
  assign acc_10_nl = { FpAdd_8U_23U_2_a_right_shift_qelse_mux_14_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12596" *) { FpAdd_8U_23U_2_a_right_shift_qelse_mux_15_nl, 1'b1 };
  assign acc_9_nl = { FpAdd_8U_23U_2_a_right_shift_qelse_mux_12_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12603" *) { FpAdd_8U_23U_2_a_right_shift_qelse_mux_13_nl, 1'b1 };
  assign acc_5_nl = { FpAdd_8U_23U_2_a_right_shift_qelse_mux_8_nl, 1'b1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12610" *) { FpAdd_8U_23U_2_a_right_shift_qelse_mux_9_nl, 1'b1 };
  assign z_out_4 = FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13225" *) 9'b110000001;
  assign z_out_5 = FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13227" *) 9'b110000001;
  assign z_out_6 = FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13229" *) 9'b110000001;
  assign z_out_7 = FpAdd_8U_23U_o_expo_lpi_1_dfm_7 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13231" *) 9'b110000001;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s[8:0] = lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[8:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4234" *) 6'b100011;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s = lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[8:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4243" *) 6'b100011;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s[8:0] = lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[8:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4252" *) 6'b100011;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s = lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[8:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4261" *) 6'b100011;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s[8:0] = lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[8:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4270" *) 6'b100011;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s = lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[8:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4279" *) 6'b100011;
  assign { _02030_[8], nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s } = lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[8:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4288" *) 6'b100011;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s = lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[8:0] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4297" *) 6'b100011;
  assign { _02029_[7:4], lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl } = { 1'b1, _02310_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4448" *) 4'b1101;
  assign lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl = { 1'b1, _02311_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4459" *) 4'b1101;
  assign lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl = { 1'b1, _02312_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4494" *) 4'b1101;
  assign lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl = { 1'b1, _02313_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4505" *) 4'b1101;
  assign lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl = { 1'b1, _02314_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4540" *) 4'b1101;
  assign lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl = { 1'b1, _02315_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4551" *) 4'b1101;
  assign lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl = { 1'b1, _02316_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4586" *) 4'b1101;
  assign lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl = { 1'b1, _02317_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4597" *) 4'b1101;
  assign _00886_ = { reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5543" *) { 2'b11, _02331_ };
  assign lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt = _00886_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5543" *) 1'b1;
  assign lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt = { reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5546" *) 1'b1;
  assign _00887_ = { reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5593" *) { 2'b11, _02338_ };
  assign lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt = _00887_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5593" *) 1'b1;
  assign lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt = { reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5596" *) 1'b1;
  assign _00888_ = { reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5633" *) { 2'b11, _02345_ };
  assign lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt = _00888_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5633" *) 1'b1;
  assign lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt = { reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5636" *) 1'b1;
  assign _00889_ = { reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5664" *) { 2'b11, _02350_ };
  assign lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt = _00889_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5664" *) 1'b1;
  assign lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt = { reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5667" *) 1'b1;
  assign lut_lookup_1_IntLog2_32U_acc_1_nl = lut_lookup_1_IntLog2_32U_lshift_itm + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5952" *) 31'b1111111111111111111111111111111;
  assign lut_lookup_1_if_else_else_else_else_else_acc_nl = { 2'b11, nl_lut_lookup_1_IntLog2_32U_lshift_rg_s[4:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5969" *) 7'b1011101;
  assign lut_lookup_1_if_else_else_else_else_if_acc_nl = { 1'b1, reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[4:2] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5972" *) 4'b1001;
  assign lut_lookup_1_else_1_else_else_acc_nl = { cfg_lut_lo_index_select_1_sva_6[7], cfg_lut_lo_index_select_1_sva_6 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6002" *) 9'b111011101;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl = { _00066_[7], _00066_[7], _00066_[5:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6005" *) 8'b11110101;
  assign lut_lookup_2_IntLog2_32U_acc_1_nl = lut_lookup_2_IntLog2_32U_lshift_itm + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6016" *) 31'b1111111111111111111111111111111;
  assign lut_lookup_2_if_else_else_else_else_else_acc_nl = { 2'b11, nl_lut_lookup_2_IntLog2_32U_lshift_rg_s[4:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6027" *) 7'b1011101;
  assign lut_lookup_2_if_else_else_else_else_if_acc_nl = { 1'b1, reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[4:2] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6030" *) 4'b1001;
  assign lut_lookup_3_IntLog2_32U_acc_1_nl = lut_lookup_3_IntLog2_32U_lshift_itm + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6062" *) 31'b1111111111111111111111111111111;
  assign lut_lookup_3_if_else_else_else_else_else_acc_nl = { 2'b11, nl_lut_lookup_3_IntLog2_32U_lshift_rg_s[4:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6072" *) 7'b1011101;
  assign lut_lookup_3_if_else_else_else_else_if_acc_nl = { 1'b1, reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[4:2] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6075" *) 4'b1001;
  assign lut_lookup_4_IntLog2_32U_acc_1_nl = lut_lookup_4_IntLog2_32U_lshift_itm + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6104" *) 31'b1111111111111111111111111111111;
  assign lut_lookup_4_if_else_else_else_else_else_acc_nl = { 2'b11, nl_lut_lookup_4_IntLog2_32U_lshift_rg_s[4:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6114" *) 7'b1011101;
  assign lut_lookup_4_if_else_else_else_else_if_acc_nl = { 1'b1, reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[4:2] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6117" *) 4'b1001;
  assign lut_lookup_1_else_else_else_if_acc_nl = IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_1_sva[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6212" *) 4'b1111;
  assign lut_lookup_2_else_else_else_if_acc_nl = IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_2_sva[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6252" *) 4'b1111;
  assign lut_lookup_3_else_else_else_if_acc_nl = IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_3_sva[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6292" *) 4'b1111;
  assign lut_lookup_4_else_else_else_if_acc_nl = IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_sva[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6332" *) 4'b1111;
  assign lut_lookup_1_if_else_else_else_else_acc_nl = { reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], nl_lut_lookup_1_IntLog2_32U_lshift_rg_s[4:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6354" *) 33'b111111111111111111111111111011101;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0 = { _00067_[7], _00067_[7], _00067_[5:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6360" *) 8'b11110101;
  assign lut_lookup_1_if_else_else_else_if_acc_nl = { reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm, reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6364" *) 4'b1111;
  assign lut_lookup_2_if_else_else_else_else_acc_nl = { reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], nl_lut_lookup_2_IntLog2_32U_lshift_rg_s[4:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6370" *) 33'b111111111111111111111111111011101;
  assign lut_lookup_2_if_else_else_else_if_acc_nl = { reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm, reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6377" *) 4'b1111;
  assign lut_lookup_3_if_else_else_else_else_acc_nl = { reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], nl_lut_lookup_3_IntLog2_32U_lshift_rg_s[4:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6385" *) 33'b111111111111111111111111111011101;
  assign lut_lookup_3_if_else_else_else_if_acc_nl = { reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm, reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6392" *) 4'b1111;
  assign lut_lookup_4_if_else_else_else_else_acc_nl = { reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], nl_lut_lookup_4_IntLog2_32U_lshift_rg_s[4:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6400" *) 33'b111111111111111111111111111011101;
  assign lut_lookup_4_if_else_else_else_if_acc_nl = { reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm, reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6407" *) 4'b1111;
  assign lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl = lut_lookup_1_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6491" *) FpMantRNE_49U_24U_1_else_carry_1_sva_2;
  assign lut_lookup_1_else_else_else_else_acc_itm_mx0w0 = { cfg_lut_le_index_select_1_sva_6[7], cfg_lut_le_index_select_1_sva_6 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6498" *) 9'b111011101;
  assign lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl = lut_lookup_1_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6501" *) FpMantRNE_49U_24U_2_else_carry_1_sva_2;
  assign lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl = lut_lookup_2_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6508" *) FpMantRNE_49U_24U_1_else_carry_2_sva_2;
  assign lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl = lut_lookup_2_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6515" *) FpMantRNE_49U_24U_2_else_carry_2_sva_2;
  assign lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl = lut_lookup_3_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6522" *) FpMantRNE_49U_24U_1_else_carry_3_sva_2;
  assign lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl = lut_lookup_3_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6529" *) FpMantRNE_49U_24U_2_else_carry_3_sva_2;
  assign lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl = lut_lookup_4_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6536" *) FpMantRNE_49U_24U_1_else_carry_sva_2;
  assign lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl = lut_lookup_4_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6543" *) FpMantRNE_49U_24U_2_else_carry_sva_2;
  assign _00890_ = { 1'b1, cfg_lut_lo_start_rsci_d[30:23] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6555" *) _00040_;
  assign FpAdd_8U_23U_2_is_a_greater_acc_nl = _00890_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6555" *) 1'b1;
  assign _00891_ = { 1'b1, cfg_lut_lo_start_rsci_d[30:23] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6559" *) _00042_;
  assign FpAdd_8U_23U_2_is_a_greater_acc_1_nl = _00891_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6559" *) 1'b1;
  assign _00892_ = { 1'b1, cfg_lut_lo_start_rsci_d[30:23] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6563" *) _00044_;
  assign FpAdd_8U_23U_2_is_a_greater_acc_2_nl = _00892_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6563" *) 1'b1;
  assign _00893_ = { 1'b1, cfg_lut_lo_start_rsci_d[30:23] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6567" *) _00045_;
  assign FpAdd_8U_23U_2_is_a_greater_acc_3_nl = _00893_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6567" *) 1'b1;
  assign lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl = { 1'b1, FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6571" *) 1'b1;
  assign lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl = { 1'b1, FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6575" *) 1'b1;
  assign lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl = { 1'b1, FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6579" *) 1'b1;
  assign lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl = { 1'b1, FpAdd_8U_23U_2_qr_lpi_1_dfm_5[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6583" *) 1'b1;
  assign lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl = { reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6593" *) 1'b1;
  assign lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl = { 1'b1, FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6611" *) 1'b1;
  assign lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl = FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6621" *) 1'b1;
  assign lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl = { reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6644" *) 1'b1;
  assign lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl = { 1'b1, FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6664" *) 1'b1;
  assign lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl = FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6674" *) 1'b1;
  assign lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl = { reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6697" *) 1'b1;
  assign lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl = { 1'b1, FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6715" *) 1'b1;
  assign lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl = FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6725" *) 1'b1;
  assign lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl = { reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6748" *) 1'b1;
  assign lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl = { 1'b1, FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12[7:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6766" *) 1'b1;
  assign lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl = FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6776" *) 1'b1;
  assign lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = { reg_lut_lookup_1_else_else_else_else_acc_1_reg, reg_lut_lookup_1_else_else_else_else_acc_1_reg, reg_lut_lookup_1_else_else_else_else_acc_2_reg, reg_lut_lookup_1_else_else_else_else_acc_3_reg, FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_1_0_1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6799" *) { lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2[7], lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2[7], lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 };
  assign lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = { reg_lut_lookup_1_else_1_else_else_acc_1_itm[7], reg_lut_lookup_1_else_1_else_else_acc_1_itm, FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_itm_1_0_1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6802" *) { lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7], lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7], lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 };
  assign lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = { reg_lut_lookup_2_else_else_else_else_acc_1_reg, reg_lut_lookup_2_else_else_else_else_acc_1_reg, reg_lut_lookup_2_else_else_else_else_acc_2_reg, reg_lut_lookup_2_else_else_else_else_acc_3_reg, FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_2_itm_1_0_1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6811" *) { lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2[7], lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2[7], lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 };
  assign lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = { reg_lut_lookup_2_else_1_else_else_acc_1_itm[7], reg_lut_lookup_2_else_1_else_else_acc_1_itm, FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_2_itm_1_0_1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6814" *) { lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7], lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7], lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 };
  assign lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = { reg_lut_lookup_3_else_else_else_else_acc_1_reg, reg_lut_lookup_3_else_else_else_else_acc_1_reg, reg_lut_lookup_3_else_else_else_else_acc_2_reg, reg_lut_lookup_3_else_else_else_else_acc_3_reg, FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_3_itm_1_0_1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6823" *) { lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2[7], lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2[7], lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 };
  assign lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = { reg_lut_lookup_3_else_1_else_else_acc_1_itm[7], reg_lut_lookup_3_else_1_else_else_acc_1_itm, FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_3_itm_1_0_1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6826" *) { lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7], lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7], lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 };
  assign lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp = { reg_lut_lookup_4_else_else_else_else_acc_1_reg, reg_lut_lookup_4_else_else_else_else_acc_1_reg, reg_lut_lookup_4_else_else_else_else_acc_2_reg, reg_lut_lookup_4_else_else_else_else_acc_3_reg, FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_4_itm_1_0_1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6835" *) { lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2[7], lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2[7], lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 };
  assign lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp = { reg_lut_lookup_4_else_1_else_else_acc_1_itm[7], reg_lut_lookup_4_else_1_else_else_acc_1_itm, FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_4_itm_1_0_1 } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6838" *) { lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7], lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2[7], lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 };
  assign lut_lookup_1_else_if_else_if_acc_nl = lut_lookup_else_if_else_le_int_1_lpi_1_dfm_1[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6841" *) 4'b1111;
  assign lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = { 1'b1, _02441_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6874" *) 1'b1;
  assign lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = { 1'b1, _02442_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6881" *) 1'b1;
  assign lut_lookup_2_else_if_else_if_acc_nl = lut_lookup_else_if_else_le_int_2_lpi_1_dfm_1[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6899" *) 4'b1111;
  assign lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = { 1'b1, _02443_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6932" *) 1'b1;
  assign lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = { 1'b1, _02444_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6939" *) 1'b1;
  assign lut_lookup_3_else_if_else_if_acc_nl = lut_lookup_else_if_else_le_int_3_lpi_1_dfm_1[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6957" *) 4'b1111;
  assign lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = { 1'b1, _02445_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6990" *) 1'b1;
  assign lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = { 1'b1, _02446_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6997" *) 1'b1;
  assign lut_lookup_4_else_if_else_if_acc_nl = lut_lookup_else_if_else_le_int_lpi_1_dfm_1[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7015" *) 4'b1111;
  assign lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl = { 1'b1, _02447_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7048" *) 1'b1;
  assign lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl = { 1'b1, _02028_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7055" *) 1'b1;
  assign lut_lookup_1_if_if_else_else_if_acc_nl = lut_lookup_if_if_else_else_le_index_s_1_sva[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7286" *) 4'b1111;
  assign lut_lookup_2_if_if_else_else_if_acc_nl = lut_lookup_if_if_else_else_le_index_s_2_sva[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7294" *) 4'b1111;
  assign lut_lookup_3_if_if_else_else_if_acc_nl = lut_lookup_if_if_else_else_le_index_s_3_sva[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7302" *) 4'b1111;
  assign lut_lookup_4_if_if_else_else_if_acc_nl = lut_lookup_if_if_else_else_le_index_s_sva[8:6] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7310" *) 4'b1111;
  assign _00894_ = { 1'b1, cfg_lut_le_start_rsci_d[30:23] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7338" *) _00040_;
  assign FpAdd_8U_23U_1_is_a_greater_acc_4_nl = _00894_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7338" *) 1'b1;
  assign _00895_ = { 1'b1, cfg_lut_le_start_rsci_d[30:23] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7342" *) _00042_;
  assign FpAdd_8U_23U_1_is_a_greater_acc_6_nl = _00895_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7342" *) 1'b1;
  assign _00896_ = { 1'b1, cfg_lut_le_start_rsci_d[30:23] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7346" *) _00044_;
  assign FpAdd_8U_23U_1_is_a_greater_acc_8_nl = _00896_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7346" *) 1'b1;
  assign _00897_ = { 1'b1, cfg_lut_le_start_rsci_d[30:23] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7350" *) _00045_;
  assign FpAdd_8U_23U_1_is_a_greater_acc_10_nl = _00897_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7350" *) 1'b1;
  assign _00898_ = { 1'b1, chn_lut_in_rsci_d_mxwt[22:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7354" *) _00068_;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl = _00898_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7354" *) 1'b1;
  assign _00899_ = { 1'b1, chn_lut_in_rsci_d_mxwt[54:32] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7358" *) _00068_;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl = _00899_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7358" *) 1'b1;
  assign _00900_ = { 1'b1, chn_lut_in_rsci_d_mxwt[86:64] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7362" *) _00068_;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl = _00900_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7362" *) 1'b1;
  assign _00901_ = { 1'b1, chn_lut_in_rsci_d_mxwt[118:96] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7366" *) _00068_;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl = _00901_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7366" *) 1'b1;
  assign lut_lookup_1_else_else_else_else_le_data_f_acc_2 = lut_lookup_1_else_else_else_else_le_data_f_lshift_1_itm + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7370" *) 32'd4294967295;
  assign lut_lookup_1_else_1_else_else_lo_data_f_acc_2 = lut_lookup_1_else_1_else_else_lo_data_f_lshift_1_itm + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7373" *) 32'd4294967295;
  assign _00902_ = { 1'b1, _02465_, _02466_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7377" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12;
  assign lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl = _00902_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7377" *) 1'b1;
  assign _00903_ = { 1'b1, _02467_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7383" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13;
  assign lut_lookup_1_FpNormalize_8U_49U_2_acc_nl = _00903_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7383" *) 1'b1;
  assign _00904_ = { 1'b1, _02468_, _02469_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7389" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14;
  assign lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl = _00904_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7389" *) 1'b1;
  assign _00905_ = { 1'b1, _02470_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7395" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15;
  assign lut_lookup_2_FpNormalize_8U_49U_2_acc_nl = _00905_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7395" *) 1'b1;
  assign _00906_ = { 1'b1, _02471_, _02472_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7401" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_16;
  assign lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl = _00906_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7401" *) 1'b1;
  assign _00907_ = { 1'b1, _02473_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7407" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_17;
  assign lut_lookup_3_FpNormalize_8U_49U_2_acc_nl = _00907_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7407" *) 1'b1;
  assign _00908_ = { 1'b1, _02474_, _02475_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7413" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_18;
  assign lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl = _00908_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7413" *) 1'b1;
  assign _00909_ = { 1'b1, _02476_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7419" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_19;
  assign lut_lookup_4_FpNormalize_8U_49U_2_acc_nl = _00909_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7419" *) 1'b1;
  assign lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl = { 1'b1, reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7424" *) 1'b1;
  assign lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl = { 1'b1, reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7428" *) 1'b1;
  assign lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl = { 1'b1, reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7432" *) 1'b1;
  assign lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl = { 1'b1, reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm, reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7436" *) 1'b1;
  assign lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl = { 1'b1, reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7440" *) 1'b1;
  assign lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl = { 1'b1, reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7444" *) 1'b1;
  assign lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl = { 1'b1, reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7448" *) 1'b1;
  assign lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl = { 1'b1, reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5:1] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7452" *) 1'b1;
  assign _00910_ = { 1'b1, chn_lut_in_rsci_d_mxwt[22:0] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7774" *) _00069_;
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl = _00910_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7774" *) 1'b1;
  assign _00911_ = { 1'b1, chn_lut_in_rsci_d_mxwt[54:32] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7778" *) _00069_;
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl = _00911_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7778" *) 1'b1;
  assign _00912_ = { 1'b1, chn_lut_in_rsci_d_mxwt[86:64] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7782" *) _00069_;
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl = _00912_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7782" *) 1'b1;
  assign _00913_ = { 1'b1, chn_lut_in_rsci_d_mxwt[118:96] } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7786" *) _00069_;
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl = _00913_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7786" *) 1'b1;
  assign lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = { 1'b1, _02520_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7790" *) 4'b1101;
  assign lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = { 1'b1, _02521_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7793" *) 4'b1101;
  assign lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = { 1'b1, _02522_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7796" *) 4'b1101;
  assign lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = { 1'b1, _02523_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7799" *) 4'b1101;
  assign lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = { 1'b1, _02524_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7802" *) 4'b1101;
  assign lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = { 1'b1, _02525_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7805" *) 4'b1101;
  assign lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1 = { 1'b1, _02526_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7808" *) 4'b1101;
  assign lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1 = { 1'b1, _02527_ } + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7811" *) 4'b1101;
  assign _00914_ = lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10013" *) lut_lookup_else_1_slc_32_mdf_sva_8;
  assign _00915_ = lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10016" *) lut_lookup_else_1_slc_32_mdf_3_sva_8;
  assign _00916_ = lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10047" *) lut_lookup_else_1_slc_32_mdf_2_sva_8;
  assign _00917_ = lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10050" *) lut_lookup_else_1_slc_32_mdf_1_sva_8;
  assign _00918_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10057" *) lut_lookup_else_else_lut_lookup_else_else_or_3_cse;
  assign _00919_ = _00918_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10058" *) mux_372_nl;
  assign _00920_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10108" *) lut_lookup_FpAdd_8U_23U_2_or_9_cse;
  assign _00921_ = _00920_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10108" *) _02100_;
  assign _00922_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10117" *) lut_lookup_FpAdd_8U_23U_2_or_8_cse;
  assign _00923_ = _00922_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10117" *) _02100_;
  assign _00925_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10204" *) _02102_;
  assign _00926_ = _00920_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10212" *) _02102_;
  assign _00927_ = _00922_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10230" *) _02103_;
  assign _00928_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10282" *) IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_5_cse;
  assign _00929_ = _00928_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10283" *) not_tmp_47;
  assign _00930_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10308" *) _02619_;
  assign _00931_ = _00930_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10308" *) not_tmp_47;
  assign _00932_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10319" *) _02622_;
  assign _00933_ = _00932_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10319" *) _02105_;
  assign _00934_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10330" *) _02624_;
  assign _00935_ = _00934_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10330" *) _02107_;
  assign _00936_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10341" *) _02627_;
  assign _00937_ = _00936_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10341" *) _02108_;
  assign _00938_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10352" *) _02629_;
  assign _00939_ = _00938_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10352" *) _02107_;
  assign _00940_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10363" *) _02632_;
  assign _00941_ = _00940_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10363" *) _02109_;
  assign _00942_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10374" *) _02634_;
  assign _00943_ = _00942_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10374" *) _02107_;
  assign _00944_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10385" *) _02637_;
  assign _00945_ = _00944_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10385" *) _02110_;
  assign _00946_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10395" *) mux_653_nl;
  assign _00947_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10403" *) mux_654_nl;
  assign _00948_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10411" *) mux_655_nl;
  assign _00949_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10419" *) mux_657_nl;
  assign _00950_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10427" *) mux_658_nl;
  assign _00951_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10435" *) mux_659_nl;
  assign _00952_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10443" *) mux_660_nl;
  assign _00953_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10451" *) mux_661_nl;
  assign _00954_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10459" *) IsNaN_8U_23U_5_IsNaN_8U_23U_6_aelse_or_2_cse;
  assign _00955_ = _00954_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10460" *) mux_667_nl;
  assign _00956_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10483" *) mux_672_nl;
  assign _00957_ = _00954_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10492" *) mux_678_nl;
  assign _00958_ = _00954_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10504" *) mux_689_nl;
  assign _00959_ = _00954_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10516" *) mux_700_nl;
  assign _00960_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10526" *) _02111_;
  assign _00962_ = _00961_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10553" *) mux_711_nl;
  assign _00963_ = _00961_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10573" *) mux_722_nl;
  assign _00964_ = _00961_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10601" *) mux_732_nl;
  assign _00965_ = _00961_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10621" *) mux_739_nl;
  assign _00966_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10642" *) mux_759_nl;
  assign _00967_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10650" *) mux_768_nl;
  assign _00968_ = and_dcpl_648 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10670" *) _02112_;
  assign _00969_ = _00968_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10670" *) or_1857_cse;
  assign _00970_ = _00969_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10671" *) lut_lookup_1_if_else_slc_32_svs_7;
  assign _00971_ = _00970_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10672" *) _02113_;
  assign _00972_ = _00971_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10672" *) FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6;
  assign _00973_ = _00972_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10673" *) lut_lookup_1_if_else_else_else_if_acc_nl[3];
  assign _00974_ = _00973_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10673" *) _02114_;
  assign _00975_ = mux_1246_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10681" *) and_dcpl_648;
  assign _00976_ = _00975_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10681" *) or_cse;
  assign _00977_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10690" *) mux_783_nl;
  assign _00978_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10699" *) mux_784_nl;
  assign _00979_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10707" *) mux_785_nl;
  assign _00980_ = lut_lookup_else_else_else_le_index_u_1_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10709" *) lut_lookup_1_else_else_else_else_le_data_f_acc_2;
  assign _00981_ = _02640_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10745" *) or_cse;
  assign _00982_ = _00981_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10745" *) core_wen;
  assign _00983_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10773" *) mux_792_nl;
  assign _00984_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10781" *) mux_797_nl;
  assign _00985_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10789" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_7;
  assign _00986_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10790" *) _02641_;
  assign _00987_ = _00986_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10790" *) _02116_;
  assign _00988_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10799" *) _02117_;
  assign _00989_ = lut_lookup_else_1_lo_index_u_1_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10801" *) lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
  assign _00990_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10808" *) _02118_;
  assign _00991_ = _00990_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10808" *) main_stage_v_3;
  assign _00992_ = _00991_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10809" *) or_1857_cse;
  assign _00993_ = _00992_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10809" *) lut_lookup_else_1_slc_32_mdf_1_sva_7;
  assign _00994_ = _00993_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10810" *) _02119_;
  assign _00995_ = _00994_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10810" *) FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5;
  assign _00996_ = _00995_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10810" *) or_cse;
  assign _00997_ = _02120_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10818" *) core_wen;
  assign _00998_ = _00997_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10818" *) _02118_;
  assign _00999_ = _00998_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10819" *) main_stage_v_3;
  assign _01000_ = _00999_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10819" *) or_cse;
  assign _01001_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10828" *) mux_803_nl;
  assign _01002_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10837" *) mux_806_nl;
  assign _01003_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10845" *) mux_823_nl;
  assign _01004_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10853" *) mux_832_nl;
  assign _01005_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10874" *) mux_840_nl;
  assign _01006_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10883" *) mux_841_nl;
  assign { _02027_[31:6], _01007_ } = lut_lookup_else_else_else_le_index_u_2_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10885" *) lut_lookup_1_else_else_else_else_le_data_f_acc_2;
  assign _01008_ = _02642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10893" *) or_cse;
  assign _01009_ = _01008_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10893" *) core_wen;
  assign _01010_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10901" *) mux_848_nl;
  assign _01011_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10921" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_7;
  assign _01012_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10922" *) _02643_;
  assign _01013_ = _01012_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10922" *) _02122_;
  assign _01014_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10931" *) _02123_;
  assign _01015_ = lut_lookup_else_1_lo_index_u_2_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10933" *) lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
  assign _01016_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10940" *) _02124_;
  assign _01017_ = _01016_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10940" *) main_stage_v_3;
  assign _01018_ = _01017_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10941" *) or_1857_cse;
  assign _01019_ = _01018_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10941" *) lut_lookup_else_1_slc_32_mdf_2_sva_7;
  assign _01020_ = _01019_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10942" *) _02125_;
  assign _01021_ = _01020_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10942" *) FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5;
  assign _01022_ = _01021_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10942" *) or_cse;
  assign _01023_ = _02126_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10950" *) core_wen;
  assign _01024_ = _01023_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10950" *) _02124_;
  assign _01025_ = _01024_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10951" *) main_stage_v_3;
  assign _01026_ = _01025_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10951" *) or_cse;
  assign _01027_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10960" *) mux_859_nl;
  assign _01028_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10969" *) mux_861_nl;
  assign _01029_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10977" *) mux_878_nl;
  assign _01030_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10985" *) mux_887_nl;
  assign _01031_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10994" *) mux_895_nl;
  assign _01032_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11003" *) mux_896_nl;
  assign _01033_ = lut_lookup_else_else_else_le_index_u_3_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11005" *) lut_lookup_1_else_else_else_else_le_data_f_acc_2;
  assign _01034_ = _02644_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11013" *) or_cse;
  assign _01035_ = _01034_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11013" *) core_wen;
  assign _01036_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11021" *) mux_903_nl;
  assign _01037_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11029" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_7;
  assign _01038_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11030" *) _02645_;
  assign _01039_ = _01038_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11030" *) _02128_;
  assign _01040_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11039" *) _02129_;
  assign _01041_ = lut_lookup_else_1_lo_index_u_3_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11041" *) lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
  assign _01042_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11048" *) _02130_;
  assign _01043_ = _01042_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11048" *) main_stage_v_3;
  assign _01044_ = _01043_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11049" *) or_1857_cse;
  assign _01045_ = _01044_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11049" *) lut_lookup_else_1_slc_32_mdf_3_sva_7;
  assign _01046_ = _01045_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11050" *) _02131_;
  assign _01047_ = _01046_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11050" *) FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5;
  assign _01048_ = _01047_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11050" *) or_cse;
  assign _01049_ = mux_1251_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11058" *) core_wen;
  assign _01050_ = _01049_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11058" *) _02130_;
  assign _01051_ = _01050_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11059" *) main_stage_v_3;
  assign _01052_ = _01051_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11059" *) or_cse;
  assign _01053_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11068" *) mux_916_nl;
  assign _01054_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11087" *) mux_926_nl;
  assign _01055_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11095" *) mux_936_nl;
  assign _01056_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11103" *) mux_945_nl;
  assign _01057_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11111" *) mux_953_nl;
  assign _01058_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11120" *) mux_954_nl;
  assign _01059_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11129" *) mux_955_nl;
  assign _01060_ = lut_lookup_else_else_else_le_index_u_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11131" *) lut_lookup_1_else_else_else_else_le_data_f_acc_2;
  assign _01061_ = _02646_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11139" *) or_cse;
  assign _01062_ = _01061_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11139" *) core_wen;
  assign _01063_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11147" *) mux_962_nl;
  assign _01064_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11155" *) IsNaN_8U_23U_7_land_lpi_1_dfm_7;
  assign _01065_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11156" *) _02647_;
  assign _01066_ = _01065_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11156" *) _02133_;
  assign _01067_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11165" *) _02134_;
  assign _01068_ = lut_lookup_else_1_lo_index_u_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11167" *) lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
  assign _01069_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11174" *) _02135_;
  assign _01070_ = _01069_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11174" *) main_stage_v_3;
  assign _01071_ = _01070_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11175" *) or_1857_cse;
  assign _01072_ = _01071_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11175" *) lut_lookup_else_1_slc_32_mdf_sva_7;
  assign _01073_ = _01072_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11176" *) _02136_;
  assign _01074_ = _01073_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11176" *) FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5;
  assign _01075_ = _01074_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11176" *) or_cse;
  assign _01076_ = mux_1252_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11184" *) core_wen;
  assign _01077_ = _01076_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11184" *) _02135_;
  assign _01078_ = _01077_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11185" *) main_stage_v_3;
  assign _01079_ = _01078_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11185" *) or_cse;
  assign _01080_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11194" *) mux_975_nl;
  assign _01081_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11218" *) _02648_;
  assign _01082_ = _01081_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11218" *) mux_tmp_978;
  assign _01083_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11227" *) mux_981_nl;
  assign _01084_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11235" *) mux_986_nl;
  assign _01085_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11243" *) mux_995_nl;
  assign _01086_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11251" *) mux_997_nl;
  assign _01087_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11271" *) mux_1013_nl;
  assign _01088_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11279" *) mux_1015_nl;
  assign _01089_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11287" *) mux_1031_nl;
  assign _01090_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11295" *) mux_1033_nl;
  assign _01091_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11303" *) mux_1049_nl;
  assign _01092_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11311" *) mux_1051_nl;
  assign _01093_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11329" *) mux_1055_nl;
  assign _01094_ = lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[7:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11351" *) { _02141_, _02141_, _02141_, _02141_, _02141_, _02141_, _02141_, _02141_ };
  assign _01095_ = _01094_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11351" *) { lut_lookup_else_1_slc_32_mdf_sva_6, lut_lookup_else_1_slc_32_mdf_sva_6, lut_lookup_else_1_slc_32_mdf_sva_6, lut_lookup_else_1_slc_32_mdf_sva_6, lut_lookup_else_1_slc_32_mdf_sva_6, lut_lookup_else_1_slc_32_mdf_sva_6, lut_lookup_else_1_slc_32_mdf_sva_6, lut_lookup_else_1_slc_32_mdf_sva_6 };
  assign _01096_ = lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[7:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11354" *) { _02142_, _02142_, _02142_, _02142_, _02142_, _02142_, _02142_, _02142_ };
  assign _01097_ = _01096_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11354" *) { lut_lookup_else_1_slc_32_mdf_3_sva_6, lut_lookup_else_1_slc_32_mdf_3_sva_6, lut_lookup_else_1_slc_32_mdf_3_sva_6, lut_lookup_else_1_slc_32_mdf_3_sva_6, lut_lookup_else_1_slc_32_mdf_3_sva_6, lut_lookup_else_1_slc_32_mdf_3_sva_6, lut_lookup_else_1_slc_32_mdf_3_sva_6, lut_lookup_else_1_slc_32_mdf_3_sva_6 };
  assign _01098_ = lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[7:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11357" *) { _02143_, _02143_, _02143_, _02143_, _02143_, _02143_, _02143_, _02143_ };
  assign _01099_ = _01098_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11357" *) { lut_lookup_else_1_slc_32_mdf_2_sva_6, lut_lookup_else_1_slc_32_mdf_2_sva_6, lut_lookup_else_1_slc_32_mdf_2_sva_6, lut_lookup_else_1_slc_32_mdf_2_sva_6, lut_lookup_else_1_slc_32_mdf_2_sva_6, lut_lookup_else_1_slc_32_mdf_2_sva_6, lut_lookup_else_1_slc_32_mdf_2_sva_6, lut_lookup_else_1_slc_32_mdf_2_sva_6 };
  assign _01100_ = lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[7:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11360" *) { _02144_, _02144_, _02144_, _02144_, _02144_, _02144_, _02144_, _02144_ };
  assign _01101_ = _01100_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11360" *) { lut_lookup_else_1_slc_32_mdf_1_sva_6, lut_lookup_else_1_slc_32_mdf_1_sva_6, lut_lookup_else_1_slc_32_mdf_1_sva_6, lut_lookup_else_1_slc_32_mdf_1_sva_6, lut_lookup_else_1_slc_32_mdf_1_sva_6, lut_lookup_else_1_slc_32_mdf_1_sva_6, lut_lookup_else_1_slc_32_mdf_1_sva_6, lut_lookup_else_1_slc_32_mdf_1_sva_6 };
  assign _01102_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11375" *) lut_lookup_FpAdd_8U_23U_1_or_11_cse;
  assign _01103_ = _01102_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11375" *) mux_1058_nl;
  assign _01104_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11384" *) mux_1059_nl;
  assign _01105_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11392" *) IsZero_8U_23U_1_IsZero_8U_23U_4_or_3_cse;
  assign _01106_ = _01105_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11393" *) mux_1060_nl;
  assign _01107_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11402" *) mux_1061_nl;
  assign _01108_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11411" *) mux_1062_nl;
  assign _01109_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11420" *) lut_lookup_FpAdd_8U_23U_2_or_10_cse;
  assign _01110_ = _01109_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11420" *) mux_1063_nl;
  assign _01111_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11429" *) mux_1064_nl;
  assign _01112_ = _00920_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11438" *) mux_1066_nl;
  assign _01113_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11457" *) mux_1069_nl;
  assign _01114_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11466" *) mux_1070_nl;
  assign _01115_ = _01105_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11475" *) mux_1071_nl;
  assign _01116_ = _00922_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11484" *) mux_1073_nl;
  assign _01117_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11504" *) IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_3_aelse_or_3_cse;
  assign _01118_ = _01117_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11505" *) mux_1077_nl;
  assign _01119_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11515" *) mux_1078_nl;
  assign _01120_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11523" *) _02147_;
  assign _01121_ = _01117_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11533" *) mux_1084_nl;
  assign _01122_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11543" *) mux_1085_nl;
  assign _01123_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11551" *) _02148_;
  assign _01124_ = _01117_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11561" *) mux_1091_nl;
  assign _01125_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11571" *) mux_1092_nl;
  assign _01126_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11579" *) _02149_;
  assign _01127_ = _01117_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11589" *) mux_1096_nl;
  assign _01128_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11599" *) mux_1097_nl;
  assign _01129_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11607" *) _02150_;
  assign _01130_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11615" *) _02151_;
  assign _01131_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11623" *) mux_1103_nl;
  assign _01132_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11631" *) mux_1104_nl;
  assign _01133_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11649" *) mux_1107_nl;
  assign _01134_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11657" *) mux_1110_nl;
  assign _01135_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11665" *) mux_1112_nl;
  assign _01136_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11685" *) mux_1118_nl;
  assign lut_lookup_else_2_else_lut_lookup_else_2_else_and_nl = lut_lookup_else_2_else_else_mux_61_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11718" *) lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse;
  assign lut_lookup_else_2_else_lut_lookup_else_2_else_and_2_nl = lut_lookup_else_2_else_else_mux_60_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11726" *) lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse;
  assign lut_lookup_else_2_else_lut_lookup_else_2_else_and_4_nl = lut_lookup_else_2_else_else_mux_59_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11734" *) lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse;
  assign lut_lookup_else_2_else_lut_lookup_else_2_else_and_6_nl = lut_lookup_else_2_else_else_mux_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11742" *) lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse;
  assign _01137_ = lut_lookup_else_if_else_le_int_1_lpi_1_dfm_1[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11747" *) { lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3] };
  assign lut_lookup_else_if_lut_lookup_else_if_and_2_nl = _01137_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11747" *) { _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34] };
  assign _01138_ = lut_lookup_else_if_else_le_int_2_lpi_1_dfm_1[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11750" *) { lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3] };
  assign lut_lookup_else_if_lut_lookup_else_if_and_5_nl = _01138_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11750" *) { _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34] };
  assign _01139_ = lut_lookup_else_if_else_le_int_3_lpi_1_dfm_1[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11753" *) { lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3] };
  assign lut_lookup_else_if_lut_lookup_else_if_and_8_nl = _01139_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11753" *) { _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34] };
  assign _01140_ = lut_lookup_else_if_else_le_int_lpi_1_dfm_1[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11756" *) { lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3] };
  assign lut_lookup_else_if_lut_lookup_else_if_and_11_nl = _01140_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11756" *) { _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34] };
  assign _01141_ = lut_lookup_else_2_else_else_if_mux_5_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11759" *) lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse;
  assign lut_lookup_else_2_lut_lookup_else_2_and_4_nl = _01141_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11759" *) _02152_;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_1_nl = lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11775" *) cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_3_nl = lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11777" *) lut_lookup_le_miss_1_sva;
  assign lut_lookup_if_2_lut_lookup_if_2_and_8_nl = lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11785" *) cfg_lut_uflow_priority_1_sva_10;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_nl = lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11787" *) cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_2_nl = lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11789" *) lut_lookup_le_miss_1_sva;
  assign lut_lookup_if_2_lut_lookup_if_2_and_9_nl = lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11797" *) cfg_lut_uflow_priority_1_sva_10;
  assign _01142_ = lut_lookup_else_2_else_else_if_mux_12_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11800" *) lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse;
  assign lut_lookup_else_2_lut_lookup_else_2_and_5_nl = _01142_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11800" *) _02153_;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_3_nl = lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11816" *) cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_7_nl = lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11818" *) lut_lookup_le_miss_2_sva;
  assign lut_lookup_if_2_lut_lookup_if_2_and_10_nl = lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11826" *) cfg_lut_uflow_priority_1_sva_10;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_2_nl = lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11828" *) cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_6_nl = lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11830" *) lut_lookup_le_miss_2_sva;
  assign lut_lookup_if_2_lut_lookup_if_2_and_11_nl = lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11838" *) cfg_lut_uflow_priority_1_sva_10;
  assign _01143_ = lut_lookup_else_2_else_else_if_mux_19_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11841" *) lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse;
  assign lut_lookup_else_2_lut_lookup_else_2_and_6_nl = _01143_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11841" *) _02154_;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_5_nl = lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11857" *) cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_11_nl = lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11859" *) lut_lookup_le_miss_3_sva;
  assign lut_lookup_if_2_lut_lookup_if_2_and_12_nl = lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11867" *) cfg_lut_uflow_priority_1_sva_10;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_4_nl = lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11869" *) cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_10_nl = lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11871" *) lut_lookup_le_miss_3_sva;
  assign lut_lookup_if_2_lut_lookup_if_2_and_13_nl = lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11879" *) cfg_lut_uflow_priority_1_sva_10;
  assign _01144_ = lut_lookup_else_2_else_else_if_mux_26_itm_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11882" *) lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse;
  assign lut_lookup_else_2_lut_lookup_else_2_and_7_nl = _01144_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11882" *) _02155_;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_7_nl = lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11898" *) cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_15_nl = lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11900" *) lut_lookup_le_miss_sva;
  assign lut_lookup_if_2_lut_lookup_if_2_and_14_nl = lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11908" *) cfg_lut_uflow_priority_1_sva_10;
  assign lut_lookup_else_2_if_lut_lookup_else_2_if_and_6_nl = lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11910" *) cfg_lut_oflow_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_14_nl = lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11912" *) lut_lookup_le_miss_sva;
  assign lut_lookup_if_2_lut_lookup_if_2_and_15_nl = lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11920" *) cfg_lut_uflow_priority_1_sva_10;
  assign _01145_ = reg_cfg_precision_1_sva_st_13_cse_1[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12040" *) or_1936_cse;
  assign and_868_nl = reg_cfg_lut_le_function_1_sva_st_20_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12044" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign and_869_nl = cfg_lut_le_function_1_sva_st_41 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12046" *) FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6;
  assign and_45_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12063" *) mux_65_nl;
  assign and_864_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12111" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign and_865_nl = cfg_lut_le_function_1_sva_st_41 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12113" *) FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6;
  assign and_48_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12131" *) mux_127_nl;
  assign and_49_nl = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12142" *) mux_tmp_128;
  assign _01146_ = reg_cfg_precision_1_sva_st_13_cse_1[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12170" *) or_tmp_1692;
  assign and_861_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12174" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign and_862_nl = cfg_lut_le_function_1_sva_st_41 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12176" *) FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6;
  assign and_54_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12193" *) mux_163_nl;
  assign _01147_ = reg_cfg_precision_1_sva_st_13_cse_1[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12235" *) or_tmp_1705;
  assign and_858_nl = reg_cfg_lut_le_function_1_sva_st_20_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12239" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign and_859_nl = cfg_lut_le_function_1_sva_st_41 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12241" *) FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6;
  assign and_59_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12259" *) mux_206_nl;
  assign _01148_ = lut_lookup_4_FpMantRNE_49U_24U_2_else_and_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12271" *) main_stage_v_2;
  assign _01149_ = _01148_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12271" *) and_dcpl_98;
  assign _01150_ = IsNaN_8U_23U_6_land_1_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12292" *) main_stage_v_4;
  assign and_62_nl = _01150_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12292" *) or_tmp_314;
  assign _01151_ = FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12298" *) main_stage_v_3;
  assign and_63_nl = _01151_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12298" *) or_1857_cse;
  assign _01152_ = IsNaN_8U_23U_10_land_1_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12299" *) main_stage_v_4;
  assign and_64_nl = _01152_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12299" *) or_tmp_314;
  assign _01153_ = IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12313" *) main_stage_v_4;
  assign and_69_nl = _01153_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12313" *) or_tmp_314;
  assign _01154_ = FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12319" *) or_1857_cse;
  assign and_70_nl = _01154_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12319" *) main_stage_v_3;
  assign _01155_ = IsNaN_8U_23U_10_land_2_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12320" *) main_stage_v_4;
  assign and_71_nl = _01155_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12320" *) or_tmp_314;
  assign _01156_ = IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12333" *) main_stage_v_4;
  assign and_74_nl = _01156_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12333" *) or_tmp_314;
  assign and_75_nl = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12338" *) and_tmp_6;
  assign _01157_ = IsNaN_8U_23U_10_land_3_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12339" *) main_stage_v_4;
  assign and_76_nl = _01157_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12339" *) or_tmp_314;
  assign _01158_ = IsNaN_8U_23U_6_land_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12353" *) main_stage_v_4;
  assign and_79_nl = _01158_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12353" *) or_tmp_314;
  assign and_80_nl = FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12359" *) and_tmp_6;
  assign _01159_ = IsNaN_8U_23U_10_land_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12360" *) main_stage_v_4;
  assign and_81_nl = _01159_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12360" *) or_tmp_314;
  assign _01160_ = cfg_lut_uflow_priority_1_sva_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12372" *) lut_lookup_lo_uflow_1_lpi_1_dfm_3;
  assign and_447_nl = _01160_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12372" *) mux_tmp_1130;
  assign _01161_ = cfg_lut_uflow_priority_1_sva_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12419" *) lut_lookup_lo_uflow_2_lpi_1_dfm_3;
  assign and_451_nl = _01161_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12419" *) mux_tmp_1143;
  assign _01162_ = cfg_lut_uflow_priority_1_sva_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12474" *) lut_lookup_lo_uflow_3_lpi_1_dfm_3;
  assign and_455_nl = _01162_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12474" *) mux_tmp_1156;
  assign _01163_ = cfg_lut_uflow_priority_1_sva_9 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12517" *) lut_lookup_lo_uflow_lpi_1_dfm_3;
  assign and_459_nl = _01163_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12517" *) mux_tmp_1169;
  assign lut_lookup_else_else_lut_lookup_else_else_and_10_nl = _02219_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12558" *) lut_lookup_else_else_slc_32_mdf_sva_8;
  assign lut_lookup_if_else_lut_lookup_if_else_and_11_nl = _02220_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12560" *) lut_lookup_4_if_else_slc_32_svs_8;
  assign lut_lookup_else_else_lut_lookup_else_else_and_7_nl = _02221_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12564" *) lut_lookup_else_else_slc_32_mdf_3_sva_8;
  assign lut_lookup_if_else_lut_lookup_if_else_and_12_nl = _02222_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12566" *) lut_lookup_2_if_else_slc_32_svs_8;
  assign lut_lookup_else_else_lut_lookup_else_else_and_4_nl = _02223_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12570" *) lut_lookup_else_else_slc_32_mdf_2_sva_8;
  assign lut_lookup_if_else_lut_lookup_if_else_and_13_nl = _02224_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12572" *) lut_lookup_1_if_else_slc_32_svs_8;
  assign lut_lookup_else_else_lut_lookup_else_else_and_1_nl = _02225_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12576" *) lut_lookup_else_else_slc_32_mdf_1_sva_8;
  assign lut_lookup_if_else_lut_lookup_if_else_and_14_nl = _02226_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12578" *) lut_lookup_3_if_else_slc_32_svs_8;
  assign and_830_nl = or_1853_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12581" *) main_stage_v_4;
  assign _01164_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12628" *) _02230_;
  assign _01165_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12637" *) mux_518_nl;
  assign _01166_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12643" *) _02231_;
  assign _01167_ = or_26_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12652" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign and_827_nl = _01167_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12652" *) FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5;
  assign and_98_nl = FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12657" *) mux_548_nl;
  assign _01168_ = reg_cfg_lut_le_function_1_sva_st_19_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12660" *) FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5;
  assign _01169_ = _01168_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12660" *) or_26_cse;
  assign and_100_nl = _01169_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12660" *) main_stage_v_1;
  assign _01170_ = and_864_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12662" *) main_stage_v_2;
  assign and_101_nl = _01170_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12662" *) or_66_cse;
  assign _01171_ = FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12667" *) main_stage_v_1;
  assign and_102_nl = _01171_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12667" *) or_26_cse;
  assign and_103_nl = IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12668" *) mux_tmp_655;
  assign _01172_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12671" *) FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5;
  assign _01173_ = _01172_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12671" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign and_104_nl = _01173_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12671" *) or_26_cse;
  assign _01174_ = and_861_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12673" *) main_stage_v_2;
  assign and_105_nl = _01174_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12673" *) or_66_cse;
  assign _01175_ = FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12678" *) main_stage_v_1;
  assign and_106_nl = _01175_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12678" *) or_26_cse;
  assign _01176_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12681" *) FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5;
  assign _01177_ = _01176_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12681" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign and_108_nl = _01177_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12681" *) or_26_cse;
  assign _01178_ = and_858_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12683" *) main_stage_v_2;
  assign and_109_nl = _01178_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12683" *) or_66_cse;
  assign _01179_ = FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12688" *) main_stage_v_1;
  assign and_110_nl = _01179_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12688" *) or_26_cse;
  assign _01180_ = IsNaN_8U_23U_7_land_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12689" *) main_stage_v_2;
  assign and_111_nl = _01180_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12689" *) or_66_cse;
  assign and_112_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12698" *) mux_663_nl;
  assign and_113_nl = main_stage_v_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12709" *) mux_666_nl;
  assign and_114_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12719" *) mux_674_nl;
  assign _01181_ = lut_lookup_else_if_lor_7_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12720" *) nor_634_cse;
  assign and_115_nl = main_stage_v_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12727" *) mux_677_nl;
  assign and_116_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12736" *) mux_685_nl;
  assign _01182_ = lut_lookup_else_if_lor_6_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12737" *) nor_634_cse;
  assign and_117_nl = main_stage_v_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12744" *) mux_688_nl;
  assign and_118_nl = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12752" *) mux_696_nl;
  assign _01183_ = lut_lookup_else_if_lor_5_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12754" *) _02247_;
  assign and_119_nl = main_stage_v_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12761" *) mux_699_nl;
  assign and_823_nl = _02976_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12765" *) main_stage_v_3;
  assign and_822_nl = _02979_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12769" *) main_stage_v_3;
  assign _01184_ = lut_lookup_1_if_else_slc_32_svs_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12782" *) mux_tmp_704;
  assign and_1166_nl = mux_751_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12784" *) _02112_;
  assign _01185_ = FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12792" *) lut_lookup_1_if_else_slc_32_svs_7;
  assign and_127_nl = _01185_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12792" *) mux_tmp_704;
  assign and_1164_nl = mux_761_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12794" *) _02112_;
  assign and_819_nl = lut_lookup_1_if_else_slc_32_svs_st_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12795" *) lut_lookup_1_if_else_slc_32_svs_8;
  assign _01186_ = and_819_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12815" *) main_stage_v_4;
  assign _01187_ = _01186_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12815" *) or_tmp_314;
  assign and_815_nl = _02112_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12817" *) main_stage_v_3;
  assign and_816_nl = _02201_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12818" *) main_stage_v_4;
  assign _01188_ = lut_lookup_else_else_else_asn_mdf_1_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12821" *) lut_lookup_else_else_slc_32_mdf_1_sva_8;
  assign _01189_ = _01188_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12821" *) cfg_lut_le_function_1_sva_st_42;
  assign _01190_ = _01189_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12821" *) IsNaN_8U_23U_6_land_1_lpi_1_dfm_6;
  assign _01191_ = _01190_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12822" *) lut_lookup_else_else_else_asn_mdf_1_sva_st_3;
  assign _01192_ = _01191_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12822" *) main_stage_v_4;
  assign and_131_nl = _01192_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12822" *) or_tmp_314;
  assign and_1162_nl = mux_815_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12844" *) _02112_;
  assign _01193_ = FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12852" *) lut_lookup_2_if_else_slc_32_svs_7;
  assign and_138_nl = _01193_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12852" *) mux_tmp_704;
  assign and_1160_nl = mux_825_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12854" *) _02112_;
  assign and_812_nl = lut_lookup_2_if_else_slc_32_svs_st_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12855" *) lut_lookup_2_if_else_slc_32_svs_8;
  assign _01194_ = _01193_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12862" *) main_stage_v_3;
  assign _01195_ = _01194_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12862" *) or_1857_cse;
  assign _01196_ = lut_lookup_2_if_else_slc_32_svs_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12866" *) IsNaN_8U_23U_6_land_2_lpi_1_dfm_6;
  assign _01197_ = _01196_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *) lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _01198_ = _01197_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *) lut_lookup_2_if_else_slc_32_svs_st_5;
  assign _01199_ = _01198_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *) main_stage_v_4;
  assign _01200_ = _01199_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *) or_tmp_314;
  assign _01201_ = lut_lookup_else_else_else_asn_mdf_2_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12870" *) cfg_lut_le_function_1_sva_st_42;
  assign _01202_ = _01201_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12870" *) lut_lookup_else_else_else_asn_mdf_2_sva_st_3;
  assign _01203_ = _01202_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12871" *) lut_lookup_else_else_slc_32_mdf_2_sva_8;
  assign _01204_ = _01203_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12871" *) IsNaN_8U_23U_6_land_2_lpi_1_dfm_6;
  assign _01205_ = _01204_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12871" *) main_stage_v_4;
  assign and_142_nl = _01205_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12871" *) or_tmp_314;
  assign and_1089_nl = or_1857_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12883" *) _03020_;
  assign _01206_ = _01154_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12887" *) lut_lookup_else_1_slc_32_mdf_2_sva_7;
  assign and_147_nl = _01206_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12887" *) main_stage_v_3;
  assign and_1158_nl = mux_870_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12891" *) _02112_;
  assign _01207_ = FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12899" *) lut_lookup_3_if_else_slc_32_svs_7;
  assign and_149_nl = _01207_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12899" *) mux_tmp_704;
  assign and_1156_nl = mux_880_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12901" *) _02112_;
  assign and_808_nl = lut_lookup_3_if_else_slc_32_svs_st_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12902" *) lut_lookup_3_if_else_slc_32_svs_8;
  assign _01208_ = lut_lookup_3_if_else_slc_32_svs_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12913" *) IsNaN_8U_23U_6_land_3_lpi_1_dfm_6;
  assign _01209_ = _01208_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *) lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _01210_ = _01209_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *) lut_lookup_3_if_else_slc_32_svs_st_5;
  assign _01211_ = _01210_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *) main_stage_v_4;
  assign _01212_ = _01211_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *) or_tmp_314;
  assign _01213_ = lut_lookup_else_else_else_asn_mdf_3_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12917" *) lut_lookup_else_else_else_asn_mdf_3_sva_st_3;
  assign _01214_ = _01213_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12917" *) lut_lookup_else_else_slc_32_mdf_3_sva_8;
  assign _01215_ = _01214_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12918" *) cfg_lut_le_function_1_sva_st_42;
  assign _01216_ = _01215_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12918" *) IsNaN_8U_23U_6_land_3_lpi_1_dfm_6;
  assign _01217_ = _01216_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12918" *) main_stage_v_4;
  assign and_152_nl = _01217_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12918" *) or_tmp_314;
  assign _01218_ = or_1857_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12932" *) _03038_;
  assign nor_tmp_46 = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12936" *) lut_lookup_else_1_slc_32_mdf_3_sva_7;
  assign and_158_nl = nor_tmp_46 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12936" *) and_tmp_6;
  assign _01219_ = cfg_precision_1_sva_st_71[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12939" *) main_stage_v_4;
  assign and_1176_nl = mux_1284_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12941" *) _02201_;
  assign _01220_ = lut_lookup_4_if_else_slc_32_svs_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12945" *) mux_tmp_704;
  assign and_1153_nl = mux_1271_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12947" *) _02112_;
  assign _01221_ = FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12955" *) lut_lookup_4_if_else_slc_32_svs_7;
  assign and_160_nl = _01221_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12955" *) mux_tmp_704;
  assign and_1151_nl = mux_1270_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12957" *) _02112_;
  assign and_804_nl = lut_lookup_4_if_else_slc_32_svs_st_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12958" *) lut_lookup_4_if_else_slc_32_svs_8;
  assign and_1174_nl = mux_1283_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12964" *) _02201_;
  assign _01222_ = and_804_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12974" *) main_stage_v_4;
  assign _01223_ = _01222_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12974" *) or_tmp_314;
  assign _01224_ = lut_lookup_else_else_else_asn_mdf_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12977" *) lut_lookup_else_else_slc_32_mdf_sva_8;
  assign _01225_ = _01224_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12977" *) cfg_lut_le_function_1_sva_st_42;
  assign _01226_ = _01225_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12977" *) IsNaN_8U_23U_6_land_lpi_1_dfm_6;
  assign _01227_ = _01226_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12978" *) lut_lookup_else_else_else_asn_mdf_sva_st_3;
  assign _01228_ = _01227_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12978" *) main_stage_v_4;
  assign and_163_nl = _01228_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12978" *) or_tmp_314;
  assign _01229_ = cfg_lut_le_function_1_sva_st_42 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12982" *) IsNaN_8U_23U_6_land_lpi_1_dfm_6;
  assign _01230_ = _01229_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12982" *) lut_lookup_else_else_slc_32_mdf_sva_8;
  assign and_166_nl = _01230_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12982" *) mux_949_nl;
  assign _01231_ = or_1857_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12993" *) _03061_;
  assign _01232_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12999" *) lut_lookup_1_if_else_slc_32_svs_6;
  assign _01233_ = _01232_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12999" *) or_66_cse;
  assign and_179_nl = _01232_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13010" *) mux_tmp_655;
  assign and_1147_nl = mux_1266_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13012" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _01234_ = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13016" *) lut_lookup_2_if_else_slc_32_svs_6;
  assign _01235_ = _01234_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13016" *) or_66_cse;
  assign and_193_nl = _01234_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13026" *) mux_tmp_655;
  assign and_1149_nl = mux_1268_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13028" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _01236_ = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13032" *) lut_lookup_3_if_else_slc_32_svs_6;
  assign _01237_ = _01236_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13032" *) or_66_cse;
  assign and_204_nl = _01236_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13042" *) mux_tmp_655;
  assign and_1148_nl = mux_1267_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13044" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _01238_ = IsNaN_8U_23U_1_land_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13048" *) lut_lookup_4_if_else_slc_32_svs_6;
  assign _01239_ = _01238_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13048" *) or_66_cse;
  assign and_215_nl = _01238_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13058" *) mux_tmp_655;
  assign and_1146_nl = mux_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13060" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _01240_ = cfg_lut_le_function_rsci_d & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13074" *) chn_lut_in_rsci_bawt;
  assign _01241_ = and_795_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13079" *) cfg_lut_le_function_rsci_d;
  assign _01242_ = reg_cfg_lut_le_function_1_sva_st_19_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13080" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
  assign _01243_ = _01240_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13115" *) and_dcpl_309;
  assign _01244_ = and_780_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13121" *) cfg_lut_le_function_rsci_d;
  assign _01245_ = reg_cfg_lut_le_function_1_sva_st_19_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13122" *) reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse;
  assign _01246_ = lut_lookup_1_if_else_slc_32_svs_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13132" *) main_stage_v_2;
  assign and_219_nl = _01246_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13132" *) or_66_cse;
  assign _01247_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13134" *) main_stage_v_2;
  assign _01248_ = _01247_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13134" *) or_66_cse;
  assign _01249_ = lut_lookup_else_else_slc_32_mdf_1_sva_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13136" *) main_stage_v_3;
  assign and_220_nl = _01249_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13137" *) or_1857_cse;
  assign _01250_ = lut_lookup_1_else_else_else_if_acc_nl[3] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13143" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _01251_ = _01250_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13143" *) lut_lookup_1_if_else_slc_32_svs_6;
  assign _01252_ = _01251_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13143" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign _01253_ = _01252_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13144" *) main_stage_v_2;
  assign and_221_nl = _01253_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13144" *) or_66_cse;
  assign and_222_nl = lut_lookup_2_if_else_slc_32_svs_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13151" *) mux_tmp_655;
  assign and_224_nl = lut_lookup_else_else_slc_32_mdf_2_sva_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13155" *) mux_tmp_704;
  assign _01254_ = _01234_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13159" *) lut_lookup_2_else_else_else_if_acc_nl[3];
  assign _01255_ = _01254_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13160" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _01256_ = _01255_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13160" *) main_stage_v_2;
  assign and_226_nl = _01256_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13160" *) or_66_cse;
  assign _01257_ = lut_lookup_else_1_slc_32_mdf_2_sva_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13164" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_6;
  assign _01258_ = _01257_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13164" *) mux_tmp_655;
  assign and_228_nl = lut_lookup_3_if_else_slc_32_svs_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13168" *) mux_tmp_655;
  assign and_230_nl = lut_lookup_else_else_slc_32_mdf_3_sva_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13172" *) mux_tmp_704;
  assign _01259_ = _01236_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13176" *) lut_lookup_3_else_else_else_if_acc_nl[3];
  assign _01260_ = _01259_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13177" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _01261_ = _01260_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13177" *) main_stage_v_2;
  assign and_232_nl = _01261_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13177" *) or_66_cse;
  assign _01262_ = lut_lookup_4_if_else_slc_32_svs_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13184" *) main_stage_v_2;
  assign and_233_nl = _01262_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13184" *) or_66_cse;
  assign _01263_ = IsNaN_8U_23U_1_land_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13186" *) main_stage_v_2;
  assign _01264_ = _01263_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13186" *) or_66_cse;
  assign _01265_ = lut_lookup_else_else_slc_32_mdf_sva_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13188" *) main_stage_v_3;
  assign and_235_nl = _01265_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13188" *) or_1857_cse;
  assign _01266_ = and_858_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13194" *) lut_lookup_4_else_else_else_if_acc_nl[3];
  assign _01267_ = _01266_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13195" *) lut_lookup_4_if_else_slc_32_svs_6;
  assign _01268_ = _01267_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13195" *) main_stage_v_2;
  assign and_236_nl = _01268_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13195" *) or_66_cse;
  assign _01269_ = lut_lookup_else_1_slc_32_mdf_sva_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13198" *) IsNaN_8U_23U_7_land_lpi_1_dfm_6;
  assign nor_tmp_55 = _01269_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13199" *) main_stage_v_2;
  assign _01270_ = nor_tmp_55 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13199" *) or_66_cse;
  assign _01271_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13201" *) lut_lookup_1_if_else_slc_32_svs_5;
  assign _01272_ = FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13209" *) or_26_cse;
  assign _01273_ = _01272_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13209" *) main_stage_v_1;
  assign _01274_ = _01273_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13209" *) lut_lookup_2_if_else_slc_32_svs_5;
  assign _01275_ = _01234_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13211" *) _02299_;
  assign and_774_nl = _01275_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13211" *) and_42_cse;
  assign _01276_ = or_26_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13214" *) lut_lookup_3_if_else_slc_32_svs_5;
  assign _01277_ = _01236_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13216" *) _02299_;
  assign and_773_nl = _01277_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13216" *) and_42_cse;
  assign _01278_ = or_26_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13219" *) lut_lookup_4_if_else_slc_32_svs_5;
  assign _01279_ = _01238_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13221" *) main_stage_v_2;
  assign _01280_ = _01279_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13221" *) or_66_cse;
  assign _01281_ = lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13234" *) mux_tmp_1247;
  assign _01282_ = lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13239" *) mux_tmp_1247;
  assign lut_lookup_else_2_else_else_else_and_4_nl = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13241" *) mux_1288_nl;
  assign _01283_ = lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13247" *) mux_tmp_1250;
  assign _01284_ = lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13252" *) mux_tmp_1250;
  assign lut_lookup_else_2_else_else_else_and_5_nl = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13254" *) mux_1291_nl;
  assign _01285_ = lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13260" *) mux_tmp_1253;
  assign _01286_ = lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13265" *) mux_tmp_1253;
  assign lut_lookup_else_2_else_else_else_and_6_nl = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13267" *) mux_1294_nl;
  assign lut_lookup_else_2_else_else_else_and_7_nl = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13276" *) _02309_;
  assign _01287_ = lut_lookup_1_if_else_else_acc_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) and_347_rgt;
  assign _01288_ = lut_lookup_2_if_else_else_acc_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) and_347_rgt;
  assign _01289_ = lut_lookup_3_if_else_else_acc_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) and_347_rgt;
  assign _01290_ = lut_lookup_4_if_else_else_acc_nl[10] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) and_347_rgt;
  assign _01291_ = lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) and_466_cse;
  assign _01292_ = lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) and_466_cse;
  assign _01293_ = lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_6_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) and_466_cse;
  assign _01294_ = lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) and_466_cse;
  assign _01295_ = FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) and_525_rgt;
  assign _01296_ = FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) and_525_rgt;
  assign _01297_ = _02104_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) lut_lookup_or_18_rgt;
  assign _01298_ = _02104_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) lut_lookup_and_125_rgt;
  assign _01299_ = _02104_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) lut_lookup_and_121_rgt;
  assign _01300_ = _02104_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13288" *) lut_lookup_or_16_rgt;
  assign _01301_ = IsNaN_8U_23U_4_land_1_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) and_dcpl_148;
  assign _01302_ = IsNaN_8U_23U_4_land_2_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) and_dcpl_148;
  assign _01303_ = IsNaN_8U_23U_4_land_3_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) and_dcpl_148;
  assign _01304_ = IsNaN_8U_23U_4_land_lpi_1_dfm_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) and_dcpl_148;
  assign _01305_ = lut_lookup_if_else_lut_lookup_if_else_and_11_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) and_465_cse;
  assign _01306_ = lut_lookup_if_else_lut_lookup_if_else_and_12_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) and_465_cse;
  assign _01307_ = lut_lookup_if_else_lut_lookup_if_else_and_13_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) and_465_cse;
  assign _01308_ = lut_lookup_if_else_lut_lookup_if_else_and_14_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) and_465_cse;
  assign _01309_ = IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) and_529_rgt;
  assign _01310_ = IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) and_529_rgt;
  assign _01311_ = FpAdd_8U_23U_1_mux_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) lut_lookup_or_17_rgt;
  assign _01312_ = FpAdd_8U_23U_1_mux_17_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) lut_lookup_and_124_rgt;
  assign _01313_ = FpAdd_8U_23U_1_mux_33_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) lut_lookup_and_120_rgt;
  assign _01314_ = FpAdd_8U_23U_1_mux_49_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) lut_lookup_or_rgt;
  assign _01315_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_344_rgt;
  assign _01316_ = IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_364_rgt;
  assign _01317_ = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_364_rgt;
  assign _01318_ = IsNaN_8U_23U_1_land_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_364_rgt;
  assign _01319_ = lut_lookup_else_else_lut_lookup_else_else_and_10_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_dcpl_258;
  assign _01320_ = lut_lookup_else_else_lut_lookup_else_else_and_7_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_dcpl_258;
  assign _01321_ = lut_lookup_else_else_lut_lookup_else_else_and_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_dcpl_258;
  assign _01322_ = lut_lookup_else_else_lut_lookup_else_else_and_1_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_dcpl_258;
  assign _01323_ = IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_527_rgt;
  assign _01324_ = lut_in_data_sva_154[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_551_rgt;
  assign _01325_ = lut_in_data_sva_154[63] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_566_rgt;
  assign _01326_ = lut_in_data_sva_154[95] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_576_rgt;
  assign _01327_ = lut_in_data_sva_154[127] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) and_588_rgt;
  assign _01328_ = FpMantRNE_49U_24U_2_else_carry_1_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *) and_564_rgt;
  assign _01329_ = FpMantRNE_49U_24U_2_else_carry_2_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *) and_564_rgt;
  assign _01330_ = FpMantRNE_49U_24U_2_else_carry_3_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *) and_586_rgt;
  assign _01331_ = FpMantRNE_49U_24U_2_else_carry_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *) and_586_rgt;
  assign _01332_ = lut_lookup_if_if_lor_1_lpi_1_dfm_mx0w3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *) and_dcpl_405;
  assign _01333_ = lut_lookup_if_if_lor_7_lpi_1_dfm_mx0w3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *) and_dcpl_405;
  assign _01334_ = lut_lookup_if_if_lor_6_lpi_1_dfm_mx0w3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *) and_dcpl_405;
  assign _01335_ = lut_lookup_if_if_lor_5_lpi_1_dfm_mx0w3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13302" *) and_dcpl_405;
  assign _01336_ = _02106_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) lut_lookup_and_127_rgt;
  assign _01337_ = _02106_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) lut_lookup_and_123_rgt;
  assign _01338_ = _02106_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) lut_lookup_and_119_rgt;
  assign _01339_ = _02106_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) lut_lookup_and_113_rgt;
  assign _01340_ = FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) and_dcpl_403;
  assign _01341_ = FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) and_dcpl_403;
  assign _01342_ = FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) and_dcpl_403;
  assign _01343_ = FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) and_dcpl_403;
  assign _01344_ = FpAdd_8U_23U_2_mux_1_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) lut_lookup_and_126_rgt;
  assign _01345_ = FpAdd_8U_23U_2_mux_17_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) lut_lookup_and_122_rgt;
  assign _01346_ = FpAdd_8U_23U_2_mux_33_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) lut_lookup_and_118_rgt;
  assign _01347_ = FpAdd_8U_23U_2_mux_49_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) lut_lookup_and_112_rgt;
  assign _01348_ = lut_lookup_4_if_else_else_else_else_acc_nl[32] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) and_606_rgt;
  assign _01349_ = lut_lookup_3_if_else_else_else_else_acc_nl[32] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) and_606_rgt;
  assign _01350_ = lut_lookup_2_if_else_else_else_else_acc_nl[32] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) and_606_rgt;
  assign _01351_ = lut_lookup_1_if_else_else_else_else_acc_nl[32] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) and_606_rgt;
  assign _01352_ = lut_in_data_sva_154[31] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) and_559_rgt;
  assign _01353_ = lut_in_data_sva_154[63] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) and_570_rgt;
  assign _01354_ = lut_in_data_sva_154[95] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) and_580_rgt;
  assign _01355_ = lut_in_data_sva_154[127] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) and_595_rgt;
  assign _01356_ = IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) and_604_rgt;
  assign _01357_ = IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) and_604_rgt;
  assign _01358_ = IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) and_604_rgt;
  assign _01359_ = and_1142_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) and_604_rgt;
  assign _01360_ = lut_lookup_lo_fraction_1_lpi_1_dfm_9[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13318" *) { lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse };
  assign _01361_ = lut_lookup_lo_fraction_2_lpi_1_dfm_9[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13318" *) { lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse };
  assign _01362_ = lut_lookup_lo_fraction_3_lpi_1_dfm_9[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13318" *) { lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse };
  assign _01363_ = lut_lookup_lo_fraction_lpi_1_dfm_9[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13318" *) { lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse };
  assign _01364_ = lut_lookup_lo_fraction_1_lpi_1_dfm_1[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *) { lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse };
  assign _01365_ = lut_lookup_lo_fraction_2_lpi_1_dfm_1[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *) { lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse };
  assign _01366_ = lut_lookup_lo_fraction_3_lpi_1_dfm_1[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *) { lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse };
  assign _01367_ = lut_lookup_lo_fraction_lpi_1_dfm_1[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *) { lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse };
  assign _01368_ = lut_lookup_le_fraction_1_lpi_1_dfm_21[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *) { lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse };
  assign _01369_ = lut_lookup_le_fraction_2_lpi_1_dfm_21[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *) { lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse };
  assign _01370_ = lut_lookup_le_fraction_3_lpi_1_dfm_21[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *) { lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse };
  assign _01371_ = lut_lookup_le_fraction_lpi_1_dfm_21[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *) { lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse };
  assign _01372_ = lut_lookup_le_fraction_1_lpi_1_dfm_9[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *) { lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse };
  assign _01373_ = lut_lookup_le_fraction_2_lpi_1_dfm_9[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *) { lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse };
  assign _01374_ = lut_lookup_le_fraction_3_lpi_1_dfm_9[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *) { lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse };
  assign _01375_ = lut_lookup_le_fraction_lpi_1_dfm_9[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *) { lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse };
  assign _01376_ = lut_lookup_le_fraction_1_lpi_1_dfm_22[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *) { lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse };
  assign _01377_ = lut_lookup_le_fraction_2_lpi_1_dfm_22[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *) { lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse };
  assign _01378_ = lut_lookup_le_fraction_3_lpi_1_dfm_22[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *) { lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse };
  assign _01379_ = lut_lookup_le_fraction_lpi_1_dfm_22[11:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *) { lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse };
  assign _01380_ = lut_lookup_lo_fraction_1_lpi_1_dfm_9[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13336" *) { lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse };
  assign _01381_ = lut_lookup_lo_fraction_2_lpi_1_dfm_9[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13336" *) { lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse };
  assign _01382_ = lut_lookup_lo_fraction_3_lpi_1_dfm_9[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13336" *) { lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse };
  assign _01383_ = lut_lookup_lo_fraction_lpi_1_dfm_9[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13336" *) { lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse };
  assign _01384_ = lut_lookup_lo_fraction_1_lpi_1_dfm_1[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *) { lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse };
  assign _01385_ = lut_lookup_lo_fraction_2_lpi_1_dfm_1[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *) { lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse };
  assign _01386_ = lut_lookup_lo_fraction_3_lpi_1_dfm_1[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *) { lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse };
  assign _01387_ = lut_lookup_lo_fraction_lpi_1_dfm_1[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *) { lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse };
  assign _01388_ = lut_lookup_le_fraction_1_lpi_1_dfm_21[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *) { lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse };
  assign _01389_ = lut_lookup_le_fraction_2_lpi_1_dfm_21[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *) { lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse };
  assign _01390_ = lut_lookup_le_fraction_3_lpi_1_dfm_21[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *) { lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse };
  assign _01391_ = lut_lookup_le_fraction_lpi_1_dfm_21[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *) { lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse };
  assign _01392_ = lut_lookup_le_fraction_1_lpi_1_dfm_9[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *) { lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse };
  assign _01393_ = lut_lookup_le_fraction_2_lpi_1_dfm_9[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *) { lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse };
  assign _01394_ = lut_lookup_le_fraction_3_lpi_1_dfm_9[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *) { lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse };
  assign _01395_ = lut_lookup_le_fraction_lpi_1_dfm_9[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *) { lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse };
  assign _01396_ = lut_lookup_le_fraction_1_lpi_1_dfm_22[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *) { lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse };
  assign _01397_ = lut_lookup_le_fraction_2_lpi_1_dfm_22[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *) { lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse };
  assign _01398_ = lut_lookup_le_fraction_3_lpi_1_dfm_22[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *) { lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse };
  assign _01399_ = lut_lookup_le_fraction_lpi_1_dfm_22[34:12] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *) { lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse };
  assign _01400_ = lut_lookup_le_fraction_1_lpi_1_dfm_16_34_12_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *) { lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse };
  assign _01401_ = lut_lookup_le_fraction_2_lpi_1_dfm_16_34_12_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *) { lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse };
  assign _01402_ = lut_lookup_le_fraction_3_lpi_1_dfm_16_34_12_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *) { lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse };
  assign _01403_ = lut_lookup_le_fraction_lpi_1_dfm_16_34_12_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *) { lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse };
  assign _01404_ = lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt[7:6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13352" *) { FpAdd_8U_23U_and_43_ssc, FpAdd_8U_23U_and_43_ssc };
  assign _01405_ = lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt[7:6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13352" *) { FpAdd_8U_23U_and_45_ssc, FpAdd_8U_23U_and_45_ssc };
  assign _01406_ = lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt[7:6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13352" *) { FpAdd_8U_23U_and_47_ssc, FpAdd_8U_23U_and_47_ssc };
  assign _01407_ = lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt[7:6] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13352" *) { FpAdd_8U_23U_and_49_ssc, FpAdd_8U_23U_and_49_ssc };
  assign _01408_ = reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *) { FpAdd_8U_23U_and_51_ssc, FpAdd_8U_23U_and_51_ssc };
  assign _01409_ = reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *) { FpAdd_8U_23U_and_53_ssc, FpAdd_8U_23U_and_53_ssc };
  assign _01410_ = reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *) { FpAdd_8U_23U_and_55_ssc, FpAdd_8U_23U_and_55_ssc };
  assign _01411_ = reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *) { FpAdd_8U_23U_and_57_ssc, FpAdd_8U_23U_and_57_ssc };
  assign _01412_ = FpNormalize_8U_49U_FpNormalize_8U_49U_and_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *) { FpAdd_8U_23U_o_expo_and_3_ssc, FpAdd_8U_23U_o_expo_and_3_ssc };
  assign _01413_ = FpNormalize_8U_49U_FpNormalize_8U_49U_and_2_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *) { FpAdd_8U_23U_o_expo_and_2_ssc, FpAdd_8U_23U_o_expo_and_2_ssc };
  assign _01414_ = FpNormalize_8U_49U_FpNormalize_8U_49U_and_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *) { FpAdd_8U_23U_o_expo_and_1_ssc, FpAdd_8U_23U_o_expo_and_1_ssc };
  assign _01415_ = FpNormalize_8U_49U_FpNormalize_8U_49U_and_6_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *) { FpAdd_8U_23U_o_expo_and_ssc, FpAdd_8U_23U_o_expo_and_ssc };
  assign _01416_ = lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13366" *) { and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt, and_290_rgt };
  assign _01417_ = lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13366" *) { and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt, and_306_rgt };
  assign _01418_ = lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13366" *) { and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt, and_322_rgt };
  assign _01419_ = lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13366" *) { and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt, and_336_rgt };
  assign _01420_ = lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *) { and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt, and_288_rgt };
  assign _01421_ = lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *) { and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt, and_304_rgt };
  assign _01422_ = lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *) { and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt, and_320_rgt };
  assign _01423_ = lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *) { and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt, and_334_rgt };
  assign _01424_ = lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *) { and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt, and_286_rgt };
  assign _01425_ = lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *) { and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt, and_302_rgt };
  assign _01426_ = lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *) { and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt, and_318_rgt };
  assign _01427_ = lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *) { and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt, and_332_rgt };
  assign _01428_ = lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *) { and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt, and_284_rgt };
  assign _01429_ = lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *) { and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt, and_300_rgt };
  assign _01430_ = lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *) { and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt, and_316_rgt };
  assign _01431_ = lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *) { and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt, and_330_rgt };
  assign _01432_ = lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13380" *) { FpAdd_8U_23U_and_43_ssc, FpAdd_8U_23U_and_43_ssc, FpAdd_8U_23U_and_43_ssc, FpAdd_8U_23U_and_43_ssc, FpAdd_8U_23U_and_43_ssc, FpAdd_8U_23U_and_43_ssc };
  assign _01433_ = lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13380" *) { FpAdd_8U_23U_and_45_ssc, FpAdd_8U_23U_and_45_ssc, FpAdd_8U_23U_and_45_ssc, FpAdd_8U_23U_and_45_ssc, FpAdd_8U_23U_and_45_ssc, FpAdd_8U_23U_and_45_ssc };
  assign _01434_ = lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13380" *) { FpAdd_8U_23U_and_47_ssc, FpAdd_8U_23U_and_47_ssc, FpAdd_8U_23U_and_47_ssc, FpAdd_8U_23U_and_47_ssc, FpAdd_8U_23U_and_47_ssc, FpAdd_8U_23U_and_47_ssc };
  assign _01435_ = lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13380" *) { FpAdd_8U_23U_and_49_ssc, FpAdd_8U_23U_and_49_ssc, FpAdd_8U_23U_and_49_ssc, FpAdd_8U_23U_and_49_ssc, FpAdd_8U_23U_and_49_ssc, FpAdd_8U_23U_and_49_ssc };
  assign _01436_ = reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *) { FpAdd_8U_23U_o_expo_or_3_nl, FpAdd_8U_23U_o_expo_or_3_nl, FpAdd_8U_23U_o_expo_or_3_nl, FpAdd_8U_23U_o_expo_or_3_nl, FpAdd_8U_23U_o_expo_or_3_nl, FpAdd_8U_23U_o_expo_or_3_nl };
  assign _01437_ = reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *) { FpAdd_8U_23U_o_expo_or_2_nl, FpAdd_8U_23U_o_expo_or_2_nl, FpAdd_8U_23U_o_expo_or_2_nl, FpAdd_8U_23U_o_expo_or_2_nl, FpAdd_8U_23U_o_expo_or_2_nl, FpAdd_8U_23U_o_expo_or_2_nl };
  assign _01438_ = reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *) { FpAdd_8U_23U_o_expo_or_1_nl, FpAdd_8U_23U_o_expo_or_1_nl, FpAdd_8U_23U_o_expo_or_1_nl, FpAdd_8U_23U_o_expo_or_1_nl, FpAdd_8U_23U_o_expo_or_1_nl, FpAdd_8U_23U_o_expo_or_1_nl };
  assign _01439_ = reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *) { FpAdd_8U_23U_o_expo_or_nl, FpAdd_8U_23U_o_expo_or_nl, FpAdd_8U_23U_o_expo_or_nl, FpAdd_8U_23U_o_expo_or_nl, FpAdd_8U_23U_o_expo_or_nl, FpAdd_8U_23U_o_expo_or_nl };
  assign _01440_ = FpNormalize_8U_49U_FpNormalize_8U_49U_and_11_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *) { FpAdd_8U_23U_o_expo_and_3_ssc, FpAdd_8U_23U_o_expo_and_3_ssc, FpAdd_8U_23U_o_expo_and_3_ssc, FpAdd_8U_23U_o_expo_and_3_ssc, FpAdd_8U_23U_o_expo_and_3_ssc, FpAdd_8U_23U_o_expo_and_3_ssc };
  assign _01441_ = FpNormalize_8U_49U_FpNormalize_8U_49U_and_10_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *) { FpAdd_8U_23U_o_expo_and_2_ssc, FpAdd_8U_23U_o_expo_and_2_ssc, FpAdd_8U_23U_o_expo_and_2_ssc, FpAdd_8U_23U_o_expo_and_2_ssc, FpAdd_8U_23U_o_expo_and_2_ssc, FpAdd_8U_23U_o_expo_and_2_ssc };
  assign _01442_ = FpNormalize_8U_49U_FpNormalize_8U_49U_and_9_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *) { FpAdd_8U_23U_o_expo_and_1_ssc, FpAdd_8U_23U_o_expo_and_1_ssc, FpAdd_8U_23U_o_expo_and_1_ssc, FpAdd_8U_23U_o_expo_and_1_ssc, FpAdd_8U_23U_o_expo_and_1_ssc, FpAdd_8U_23U_o_expo_and_1_ssc };
  assign _01443_ = FpNormalize_8U_49U_FpNormalize_8U_49U_and_8_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *) { FpAdd_8U_23U_o_expo_and_ssc, FpAdd_8U_23U_o_expo_and_ssc, FpAdd_8U_23U_o_expo_and_ssc, FpAdd_8U_23U_o_expo_and_ssc, FpAdd_8U_23U_o_expo_and_ssc, FpAdd_8U_23U_o_expo_and_ssc };
  assign _01444_ = lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_13[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13396" *) { lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse, lut_lookup_and_139_cse };
  assign _01445_ = lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_13[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13396" *) { lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse, lut_lookup_and_137_cse };
  assign _01446_ = lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_13[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13396" *) { lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse, lut_lookup_and_135_cse };
  assign _01447_ = lut_lookup_lo_index_0_7_0_lpi_1_dfm_13[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13396" *) { lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse, lut_lookup_and_133_cse };
  assign _01448_ = lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_1[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *) { lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse, lut_lookup_and_138_cse };
  assign _01449_ = lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_1[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *) { lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse, lut_lookup_and_136_cse };
  assign _01450_ = lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_1[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *) { lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse, lut_lookup_and_134_cse };
  assign _01451_ = lut_lookup_lo_index_0_7_0_lpi_1_dfm_1[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *) { lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse, lut_lookup_and_132_cse };
  assign _01452_ = lut_lookup_le_index_0_5_0_1_lpi_1_dfm_26 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *) { lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse, lut_lookup_and_7_cse };
  assign _01453_ = lut_lookup_le_index_0_5_0_2_lpi_1_dfm_26 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *) { lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse, lut_lookup_and_15_cse };
  assign _01454_ = lut_lookup_le_index_0_5_0_3_lpi_1_dfm_26 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *) { lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse, lut_lookup_and_23_cse };
  assign _01455_ = lut_lookup_le_index_0_5_0_lpi_1_dfm_26 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *) { lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse, lut_lookup_and_31_cse };
  assign _01456_ = lut_lookup_else_if_lut_lookup_else_if_and_2_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *) { lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse, lut_lookup_and_6_cse };
  assign _01457_ = lut_lookup_else_if_lut_lookup_else_if_and_5_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *) { lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse, lut_lookup_and_14_cse };
  assign _01458_ = lut_lookup_else_if_lut_lookup_else_if_and_8_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *) { lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse, lut_lookup_and_22_cse };
  assign _01459_ = lut_lookup_else_if_lut_lookup_else_if_and_11_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *) { lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse, lut_lookup_and_30_cse };
  assign _01460_ = lut_lookup_le_index_0_5_0_1_lpi_1_dfm_28 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *) { lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse, lut_lookup_and_5_cse };
  assign _01461_ = lut_lookup_le_index_0_5_0_2_lpi_1_dfm_28 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *) { lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse, lut_lookup_and_13_cse };
  assign _01462_ = lut_lookup_le_index_0_5_0_3_lpi_1_dfm_28 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *) { lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse, lut_lookup_and_21_cse };
  assign _01463_ = lut_lookup_le_index_0_5_0_lpi_1_dfm_28 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *) { lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse, lut_lookup_and_29_cse };
  assign _01464_ = lut_lookup_le_index_0_5_0_1_lpi_1_dfm_29 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *) { lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse, lut_lookup_lut_lookup_nor_19_cse };
  assign _01465_ = lut_lookup_le_index_0_5_0_2_lpi_1_dfm_29 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *) { lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse, lut_lookup_lut_lookup_nor_18_cse };
  assign _01466_ = lut_lookup_le_index_0_5_0_3_lpi_1_dfm_29 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *) { lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse, lut_lookup_lut_lookup_nor_17_cse };
  assign _01467_ = lut_lookup_le_index_0_5_0_lpi_1_dfm_29 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *) { lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse, lut_lookup_lut_lookup_nor_16_cse };
  assign _01468_ = lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13412" *) { FpAdd_8U_23U_2_and_5_rgt, FpAdd_8U_23U_2_and_5_rgt, FpAdd_8U_23U_2_and_5_rgt, FpAdd_8U_23U_2_and_5_rgt, FpAdd_8U_23U_2_and_5_rgt, FpAdd_8U_23U_2_and_5_rgt, FpAdd_8U_23U_2_and_5_rgt, FpAdd_8U_23U_2_and_5_rgt };
  assign _01469_ = lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13412" *) { FpAdd_8U_23U_2_and_11_rgt, FpAdd_8U_23U_2_and_11_rgt, FpAdd_8U_23U_2_and_11_rgt, FpAdd_8U_23U_2_and_11_rgt, FpAdd_8U_23U_2_and_11_rgt, FpAdd_8U_23U_2_and_11_rgt, FpAdd_8U_23U_2_and_11_rgt, FpAdd_8U_23U_2_and_11_rgt };
  assign _01470_ = lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13412" *) { FpAdd_8U_23U_2_and_17_rgt, FpAdd_8U_23U_2_and_17_rgt, FpAdd_8U_23U_2_and_17_rgt, FpAdd_8U_23U_2_and_17_rgt, FpAdd_8U_23U_2_and_17_rgt, FpAdd_8U_23U_2_and_17_rgt, FpAdd_8U_23U_2_and_17_rgt, FpAdd_8U_23U_2_and_17_rgt };
  assign _01471_ = lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13412" *) { FpAdd_8U_23U_2_and_23_rgt, FpAdd_8U_23U_2_and_23_rgt, FpAdd_8U_23U_2_and_23_rgt, FpAdd_8U_23U_2_and_23_rgt, FpAdd_8U_23U_2_and_23_rgt, FpAdd_8U_23U_2_and_23_rgt, FpAdd_8U_23U_2_and_23_rgt, FpAdd_8U_23U_2_and_23_rgt };
  assign _01472_ = FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *) { FpAdd_8U_23U_2_and_4_rgt, FpAdd_8U_23U_2_and_4_rgt, FpAdd_8U_23U_2_and_4_rgt, FpAdd_8U_23U_2_and_4_rgt, FpAdd_8U_23U_2_and_4_rgt, FpAdd_8U_23U_2_and_4_rgt, FpAdd_8U_23U_2_and_4_rgt, FpAdd_8U_23U_2_and_4_rgt };
  assign _01473_ = FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *) { FpAdd_8U_23U_2_and_10_rgt, FpAdd_8U_23U_2_and_10_rgt, FpAdd_8U_23U_2_and_10_rgt, FpAdd_8U_23U_2_and_10_rgt, FpAdd_8U_23U_2_and_10_rgt, FpAdd_8U_23U_2_and_10_rgt, FpAdd_8U_23U_2_and_10_rgt, FpAdd_8U_23U_2_and_10_rgt };
  assign _01474_ = FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *) { FpAdd_8U_23U_2_and_16_rgt, FpAdd_8U_23U_2_and_16_rgt, FpAdd_8U_23U_2_and_16_rgt, FpAdd_8U_23U_2_and_16_rgt, FpAdd_8U_23U_2_and_16_rgt, FpAdd_8U_23U_2_and_16_rgt, FpAdd_8U_23U_2_and_16_rgt, FpAdd_8U_23U_2_and_16_rgt };
  assign _01475_ = FpAdd_8U_23U_2_qr_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *) { FpAdd_8U_23U_2_and_22_rgt, FpAdd_8U_23U_2_and_22_rgt, FpAdd_8U_23U_2_and_22_rgt, FpAdd_8U_23U_2_and_22_rgt, FpAdd_8U_23U_2_and_22_rgt, FpAdd_8U_23U_2_and_22_rgt, FpAdd_8U_23U_2_and_22_rgt, FpAdd_8U_23U_2_and_22_rgt };
  assign _01476_ = FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *) { FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt };
  assign _01477_ = FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_2_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *) { FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt };
  assign _01478_ = FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_4_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *) { FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt };
  assign _01479_ = FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_6_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *) { FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt, FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt };
  assign _01480_ = lut_in_data_sva_156[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *) { IsNaN_8U_23U_3_land_1_lpi_1_dfm_6, IsNaN_8U_23U_3_land_1_lpi_1_dfm_6, IsNaN_8U_23U_3_land_1_lpi_1_dfm_6, IsNaN_8U_23U_3_land_1_lpi_1_dfm_6, IsNaN_8U_23U_3_land_1_lpi_1_dfm_6, IsNaN_8U_23U_3_land_1_lpi_1_dfm_6, IsNaN_8U_23U_3_land_1_lpi_1_dfm_6, IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 };
  assign _01481_ = lut_in_data_sva_156[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *) { IsNaN_8U_23U_7_land_1_lpi_1_dfm_7, IsNaN_8U_23U_7_land_1_lpi_1_dfm_7, IsNaN_8U_23U_7_land_1_lpi_1_dfm_7, IsNaN_8U_23U_7_land_1_lpi_1_dfm_7, IsNaN_8U_23U_7_land_1_lpi_1_dfm_7, IsNaN_8U_23U_7_land_1_lpi_1_dfm_7, IsNaN_8U_23U_7_land_1_lpi_1_dfm_7, IsNaN_8U_23U_7_land_1_lpi_1_dfm_7 };
  assign _01482_ = lut_in_data_sva_156[62:55] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *) { IsNaN_8U_23U_3_land_2_lpi_1_dfm_7, IsNaN_8U_23U_3_land_2_lpi_1_dfm_7, IsNaN_8U_23U_3_land_2_lpi_1_dfm_7, IsNaN_8U_23U_3_land_2_lpi_1_dfm_7, IsNaN_8U_23U_3_land_2_lpi_1_dfm_7, IsNaN_8U_23U_3_land_2_lpi_1_dfm_7, IsNaN_8U_23U_3_land_2_lpi_1_dfm_7, IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 };
  assign _01483_ = lut_in_data_sva_156[62:55] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *) { IsNaN_8U_23U_7_land_2_lpi_1_dfm_7, IsNaN_8U_23U_7_land_2_lpi_1_dfm_7, IsNaN_8U_23U_7_land_2_lpi_1_dfm_7, IsNaN_8U_23U_7_land_2_lpi_1_dfm_7, IsNaN_8U_23U_7_land_2_lpi_1_dfm_7, IsNaN_8U_23U_7_land_2_lpi_1_dfm_7, IsNaN_8U_23U_7_land_2_lpi_1_dfm_7, IsNaN_8U_23U_7_land_2_lpi_1_dfm_7 };
  assign _01484_ = lut_in_data_sva_156[94:87] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *) { IsNaN_8U_23U_3_land_3_lpi_1_dfm_7, IsNaN_8U_23U_3_land_3_lpi_1_dfm_7, IsNaN_8U_23U_3_land_3_lpi_1_dfm_7, IsNaN_8U_23U_3_land_3_lpi_1_dfm_7, IsNaN_8U_23U_3_land_3_lpi_1_dfm_7, IsNaN_8U_23U_3_land_3_lpi_1_dfm_7, IsNaN_8U_23U_3_land_3_lpi_1_dfm_7, IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 };
  assign _01485_ = lut_in_data_sva_156[94:87] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *) { IsNaN_8U_23U_7_land_3_lpi_1_dfm_7, IsNaN_8U_23U_7_land_3_lpi_1_dfm_7, IsNaN_8U_23U_7_land_3_lpi_1_dfm_7, IsNaN_8U_23U_7_land_3_lpi_1_dfm_7, IsNaN_8U_23U_7_land_3_lpi_1_dfm_7, IsNaN_8U_23U_7_land_3_lpi_1_dfm_7, IsNaN_8U_23U_7_land_3_lpi_1_dfm_7, IsNaN_8U_23U_7_land_3_lpi_1_dfm_7 };
  assign _01486_ = lut_in_data_sva_156[126:119] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *) { IsNaN_8U_23U_3_land_lpi_1_dfm_6, IsNaN_8U_23U_3_land_lpi_1_dfm_6, IsNaN_8U_23U_3_land_lpi_1_dfm_6, IsNaN_8U_23U_3_land_lpi_1_dfm_6, IsNaN_8U_23U_3_land_lpi_1_dfm_6, IsNaN_8U_23U_3_land_lpi_1_dfm_6, IsNaN_8U_23U_3_land_lpi_1_dfm_6, IsNaN_8U_23U_3_land_lpi_1_dfm_6 };
  assign _01487_ = lut_in_data_sva_156[126:119] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13427" *) { IsNaN_8U_23U_7_land_lpi_1_dfm_7, IsNaN_8U_23U_7_land_lpi_1_dfm_7, IsNaN_8U_23U_7_land_lpi_1_dfm_7, IsNaN_8U_23U_7_land_lpi_1_dfm_7, IsNaN_8U_23U_7_land_lpi_1_dfm_7, IsNaN_8U_23U_7_land_lpi_1_dfm_7, IsNaN_8U_23U_7_land_lpi_1_dfm_7, IsNaN_8U_23U_7_land_lpi_1_dfm_7 };
  assign _01488_ = cfg_lut_le_start_1_sva_3_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) { FpAdd_8U_23U_and_35_nl, FpAdd_8U_23U_and_35_nl, FpAdd_8U_23U_and_35_nl, FpAdd_8U_23U_and_35_nl, FpAdd_8U_23U_and_35_nl, FpAdd_8U_23U_and_35_nl, FpAdd_8U_23U_and_35_nl, FpAdd_8U_23U_and_35_nl };
  assign _01489_ = cfg_lut_lo_start_1_sva_3_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) { FpAdd_8U_23U_2_and_9_nl, FpAdd_8U_23U_2_and_9_nl, FpAdd_8U_23U_2_and_9_nl, FpAdd_8U_23U_2_and_9_nl, FpAdd_8U_23U_2_and_9_nl, FpAdd_8U_23U_2_and_9_nl, FpAdd_8U_23U_2_and_9_nl, FpAdd_8U_23U_2_and_9_nl };
  assign _01490_ = cfg_lut_le_start_1_sva_3_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) { FpAdd_8U_23U_and_37_nl, FpAdd_8U_23U_and_37_nl, FpAdd_8U_23U_and_37_nl, FpAdd_8U_23U_and_37_nl, FpAdd_8U_23U_and_37_nl, FpAdd_8U_23U_and_37_nl, FpAdd_8U_23U_and_37_nl, FpAdd_8U_23U_and_37_nl };
  assign _01491_ = cfg_lut_lo_start_1_sva_3_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) { FpAdd_8U_23U_2_and_15_nl, FpAdd_8U_23U_2_and_15_nl, FpAdd_8U_23U_2_and_15_nl, FpAdd_8U_23U_2_and_15_nl, FpAdd_8U_23U_2_and_15_nl, FpAdd_8U_23U_2_and_15_nl, FpAdd_8U_23U_2_and_15_nl, FpAdd_8U_23U_2_and_15_nl };
  assign _01492_ = cfg_lut_le_start_1_sva_3_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) { FpAdd_8U_23U_and_39_nl, FpAdd_8U_23U_and_39_nl, FpAdd_8U_23U_and_39_nl, FpAdd_8U_23U_and_39_nl, FpAdd_8U_23U_and_39_nl, FpAdd_8U_23U_and_39_nl, FpAdd_8U_23U_and_39_nl, FpAdd_8U_23U_and_39_nl };
  assign _01493_ = cfg_lut_lo_start_1_sva_3_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) { FpAdd_8U_23U_2_and_21_nl, FpAdd_8U_23U_2_and_21_nl, FpAdd_8U_23U_2_and_21_nl, FpAdd_8U_23U_2_and_21_nl, FpAdd_8U_23U_2_and_21_nl, FpAdd_8U_23U_2_and_21_nl, FpAdd_8U_23U_2_and_21_nl, FpAdd_8U_23U_2_and_21_nl };
  assign _01494_ = cfg_lut_le_start_1_sva_3_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) { FpAdd_8U_23U_and_41_nl, FpAdd_8U_23U_and_41_nl, FpAdd_8U_23U_and_41_nl, FpAdd_8U_23U_and_41_nl, FpAdd_8U_23U_and_41_nl, FpAdd_8U_23U_and_41_nl, FpAdd_8U_23U_and_41_nl, FpAdd_8U_23U_and_41_nl };
  assign _01495_ = cfg_lut_lo_start_1_sva_3_30_0_1[30:23] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) { FpAdd_8U_23U_2_and_27_nl, FpAdd_8U_23U_2_and_27_nl, FpAdd_8U_23U_2_and_27_nl, FpAdd_8U_23U_2_and_27_nl, FpAdd_8U_23U_2_and_27_nl, FpAdd_8U_23U_2_and_27_nl, FpAdd_8U_23U_2_and_27_nl, FpAdd_8U_23U_2_and_27_nl };
  assign _01496_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) { FpAdd_8U_23U_1_and_35_nl, FpAdd_8U_23U_1_and_35_nl, FpAdd_8U_23U_1_and_35_nl, FpAdd_8U_23U_1_and_35_nl, FpAdd_8U_23U_1_and_35_nl, FpAdd_8U_23U_1_and_35_nl, FpAdd_8U_23U_1_and_35_nl, FpAdd_8U_23U_1_and_35_nl };
  assign _01497_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) { FpAdd_8U_23U_2_and_28_nl, FpAdd_8U_23U_2_and_28_nl, FpAdd_8U_23U_2_and_28_nl, FpAdd_8U_23U_2_and_28_nl, FpAdd_8U_23U_2_and_28_nl, FpAdd_8U_23U_2_and_28_nl, FpAdd_8U_23U_2_and_28_nl, FpAdd_8U_23U_2_and_28_nl };
  assign _01498_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) { FpAdd_8U_23U_1_and_37_nl, FpAdd_8U_23U_1_and_37_nl, FpAdd_8U_23U_1_and_37_nl, FpAdd_8U_23U_1_and_37_nl, FpAdd_8U_23U_1_and_37_nl, FpAdd_8U_23U_1_and_37_nl, FpAdd_8U_23U_1_and_37_nl, FpAdd_8U_23U_1_and_37_nl };
  assign _01499_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) { FpAdd_8U_23U_2_and_30_nl, FpAdd_8U_23U_2_and_30_nl, FpAdd_8U_23U_2_and_30_nl, FpAdd_8U_23U_2_and_30_nl, FpAdd_8U_23U_2_and_30_nl, FpAdd_8U_23U_2_and_30_nl, FpAdd_8U_23U_2_and_30_nl, FpAdd_8U_23U_2_and_30_nl };
  assign _01500_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) { FpAdd_8U_23U_1_and_39_nl, FpAdd_8U_23U_1_and_39_nl, FpAdd_8U_23U_1_and_39_nl, FpAdd_8U_23U_1_and_39_nl, FpAdd_8U_23U_1_and_39_nl, FpAdd_8U_23U_1_and_39_nl, FpAdd_8U_23U_1_and_39_nl, FpAdd_8U_23U_1_and_39_nl };
  assign _01501_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) { FpAdd_8U_23U_2_and_32_nl, FpAdd_8U_23U_2_and_32_nl, FpAdd_8U_23U_2_and_32_nl, FpAdd_8U_23U_2_and_32_nl, FpAdd_8U_23U_2_and_32_nl, FpAdd_8U_23U_2_and_32_nl, FpAdd_8U_23U_2_and_32_nl, FpAdd_8U_23U_2_and_32_nl };
  assign _01502_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) { FpAdd_8U_23U_1_and_41_nl, FpAdd_8U_23U_1_and_41_nl, FpAdd_8U_23U_1_and_41_nl, FpAdd_8U_23U_1_and_41_nl, FpAdd_8U_23U_1_and_41_nl, FpAdd_8U_23U_1_and_41_nl, FpAdd_8U_23U_1_and_41_nl, FpAdd_8U_23U_1_and_41_nl };
  assign _01503_ = 8'b11111110 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) { FpAdd_8U_23U_2_and_34_nl, FpAdd_8U_23U_2_and_34_nl, FpAdd_8U_23U_2_and_34_nl, FpAdd_8U_23U_2_and_34_nl, FpAdd_8U_23U_2_and_34_nl, FpAdd_8U_23U_2_and_34_nl, FpAdd_8U_23U_2_and_34_nl, FpAdd_8U_23U_2_and_34_nl };
  assign _01504_ = lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) { FpAdd_8U_23U_and_61_nl, FpAdd_8U_23U_and_61_nl, FpAdd_8U_23U_and_61_nl, FpAdd_8U_23U_and_61_nl, FpAdd_8U_23U_and_61_nl, FpAdd_8U_23U_and_61_nl, FpAdd_8U_23U_and_61_nl, FpAdd_8U_23U_and_61_nl };
  assign _01505_ = lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) { FpAdd_8U_23U_2_and_6_nl, FpAdd_8U_23U_2_and_6_nl, FpAdd_8U_23U_2_and_6_nl, FpAdd_8U_23U_2_and_6_nl, FpAdd_8U_23U_2_and_6_nl, FpAdd_8U_23U_2_and_6_nl, FpAdd_8U_23U_2_and_6_nl, FpAdd_8U_23U_2_and_6_nl };
  assign _01506_ = lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) { FpAdd_8U_23U_and_65_nl, FpAdd_8U_23U_and_65_nl, FpAdd_8U_23U_and_65_nl, FpAdd_8U_23U_and_65_nl, FpAdd_8U_23U_and_65_nl, FpAdd_8U_23U_and_65_nl, FpAdd_8U_23U_and_65_nl, FpAdd_8U_23U_and_65_nl };
  assign _01507_ = lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) { FpAdd_8U_23U_2_and_13_nl, FpAdd_8U_23U_2_and_13_nl, FpAdd_8U_23U_2_and_13_nl, FpAdd_8U_23U_2_and_13_nl, FpAdd_8U_23U_2_and_13_nl, FpAdd_8U_23U_2_and_13_nl, FpAdd_8U_23U_2_and_13_nl, FpAdd_8U_23U_2_and_13_nl };
  assign _01508_ = lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) { FpAdd_8U_23U_and_69_nl, FpAdd_8U_23U_and_69_nl, FpAdd_8U_23U_and_69_nl, FpAdd_8U_23U_and_69_nl, FpAdd_8U_23U_and_69_nl, FpAdd_8U_23U_and_69_nl, FpAdd_8U_23U_and_69_nl, FpAdd_8U_23U_and_69_nl };
  assign _01509_ = lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) { FpAdd_8U_23U_2_and_19_nl, FpAdd_8U_23U_2_and_19_nl, FpAdd_8U_23U_2_and_19_nl, FpAdd_8U_23U_2_and_19_nl, FpAdd_8U_23U_2_and_19_nl, FpAdd_8U_23U_2_and_19_nl, FpAdd_8U_23U_2_and_19_nl, FpAdd_8U_23U_2_and_19_nl };
  assign _01510_ = lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) { FpAdd_8U_23U_and_73_nl, FpAdd_8U_23U_and_73_nl, FpAdd_8U_23U_and_73_nl, FpAdd_8U_23U_and_73_nl, FpAdd_8U_23U_and_73_nl, FpAdd_8U_23U_and_73_nl, FpAdd_8U_23U_and_73_nl, FpAdd_8U_23U_and_73_nl };
  assign _01511_ = lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) { FpAdd_8U_23U_2_and_25_nl, FpAdd_8U_23U_2_and_25_nl, FpAdd_8U_23U_2_and_25_nl, FpAdd_8U_23U_2_and_25_nl, FpAdd_8U_23U_2_and_25_nl, FpAdd_8U_23U_2_and_25_nl, FpAdd_8U_23U_2_and_25_nl, FpAdd_8U_23U_2_and_25_nl };
  assign _01512_ = { reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) { FpAdd_8U_23U_and_59_nl, FpAdd_8U_23U_and_59_nl, FpAdd_8U_23U_and_59_nl, FpAdd_8U_23U_and_59_nl, FpAdd_8U_23U_and_59_nl, FpAdd_8U_23U_and_59_nl, FpAdd_8U_23U_and_59_nl, FpAdd_8U_23U_and_59_nl };
  assign _01513_ = FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) { FpAdd_8U_23U_2_and_nl, FpAdd_8U_23U_2_and_nl, FpAdd_8U_23U_2_and_nl, FpAdd_8U_23U_2_and_nl, FpAdd_8U_23U_2_and_nl, FpAdd_8U_23U_2_and_nl, FpAdd_8U_23U_2_and_nl, FpAdd_8U_23U_2_and_nl };
  assign _01514_ = { reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) { FpAdd_8U_23U_and_63_nl, FpAdd_8U_23U_and_63_nl, FpAdd_8U_23U_and_63_nl, FpAdd_8U_23U_and_63_nl, FpAdd_8U_23U_and_63_nl, FpAdd_8U_23U_and_63_nl, FpAdd_8U_23U_and_63_nl, FpAdd_8U_23U_and_63_nl };
  assign _01515_ = FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) { FpAdd_8U_23U_2_and_29_nl, FpAdd_8U_23U_2_and_29_nl, FpAdd_8U_23U_2_and_29_nl, FpAdd_8U_23U_2_and_29_nl, FpAdd_8U_23U_2_and_29_nl, FpAdd_8U_23U_2_and_29_nl, FpAdd_8U_23U_2_and_29_nl, FpAdd_8U_23U_2_and_29_nl };
  assign _01516_ = { reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) { FpAdd_8U_23U_and_67_nl, FpAdd_8U_23U_and_67_nl, FpAdd_8U_23U_and_67_nl, FpAdd_8U_23U_and_67_nl, FpAdd_8U_23U_and_67_nl, FpAdd_8U_23U_and_67_nl, FpAdd_8U_23U_and_67_nl, FpAdd_8U_23U_and_67_nl };
  assign _01517_ = FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) { FpAdd_8U_23U_2_and_31_nl, FpAdd_8U_23U_2_and_31_nl, FpAdd_8U_23U_2_and_31_nl, FpAdd_8U_23U_2_and_31_nl, FpAdd_8U_23U_2_and_31_nl, FpAdd_8U_23U_2_and_31_nl, FpAdd_8U_23U_2_and_31_nl, FpAdd_8U_23U_2_and_31_nl };
  assign _01518_ = { reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm, reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) { FpAdd_8U_23U_and_71_nl, FpAdd_8U_23U_and_71_nl, FpAdd_8U_23U_and_71_nl, FpAdd_8U_23U_and_71_nl, FpAdd_8U_23U_and_71_nl, FpAdd_8U_23U_and_71_nl, FpAdd_8U_23U_and_71_nl, FpAdd_8U_23U_and_71_nl };
  assign _01519_ = FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) { FpAdd_8U_23U_2_and_33_nl, FpAdd_8U_23U_2_and_33_nl, FpAdd_8U_23U_2_and_33_nl, FpAdd_8U_23U_2_and_33_nl, FpAdd_8U_23U_2_and_33_nl, FpAdd_8U_23U_2_and_33_nl, FpAdd_8U_23U_2_and_33_nl, FpAdd_8U_23U_2_and_33_nl };
  assign _01520_ = lut_lookup_1_if_else_else_else_else_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13444" *) { mux_1190_nl, mux_1190_nl, mux_1190_nl, mux_1190_nl, mux_1190_nl, mux_1190_nl, mux_1190_nl, mux_1190_nl, mux_1190_nl };
  assign _01521_ = lut_lookup_2_if_else_else_else_else_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13444" *) { mux_1195_nl, mux_1195_nl, mux_1195_nl, mux_1195_nl, mux_1195_nl, mux_1195_nl, mux_1195_nl, mux_1195_nl, mux_1195_nl };
  assign _01522_ = lut_lookup_3_if_else_else_else_else_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13444" *) { mux_1200_nl, mux_1200_nl, mux_1200_nl, mux_1200_nl, mux_1200_nl, mux_1200_nl, mux_1200_nl, mux_1200_nl, mux_1200_nl };
  assign _01523_ = lut_lookup_4_if_else_else_else_else_if_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13444" *) { mux_1205_nl, mux_1205_nl, mux_1205_nl, mux_1205_nl, mux_1205_nl, mux_1205_nl, mux_1205_nl, mux_1205_nl, mux_1205_nl };
  assign _01524_ = lut_lookup_1_if_else_else_else_else_else_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *) { mux_1189_nl, mux_1189_nl, mux_1189_nl, mux_1189_nl, mux_1189_nl, mux_1189_nl, mux_1189_nl, mux_1189_nl, mux_1189_nl };
  assign _01525_ = lut_lookup_2_if_else_else_else_else_else_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *) { mux_1194_nl, mux_1194_nl, mux_1194_nl, mux_1194_nl, mux_1194_nl, mux_1194_nl, mux_1194_nl, mux_1194_nl, mux_1194_nl };
  assign _01526_ = lut_lookup_3_if_else_else_else_else_else_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *) { mux_1199_nl, mux_1199_nl, mux_1199_nl, mux_1199_nl, mux_1199_nl, mux_1199_nl, mux_1199_nl, mux_1199_nl, mux_1199_nl };
  assign _01527_ = lut_lookup_4_if_else_else_else_else_else_acc_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *) { mux_1204_nl, mux_1204_nl, mux_1204_nl, mux_1204_nl, mux_1204_nl, mux_1204_nl, mux_1204_nl, mux_1204_nl, mux_1204_nl };
  assign _01528_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13446" *) { mux_1188_cse, mux_1188_cse, mux_1188_cse, mux_1188_cse, mux_1188_cse, mux_1188_cse, mux_1188_cse, mux_1188_cse, mux_1188_cse };
  assign _01529_ = z_out_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *) { and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405 };
  assign _01530_ = z_out_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *) { and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405 };
  assign _01531_ = z_out_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *) { and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405 };
  assign _01532_ = z_out_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *) { and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405, and_dcpl_405 };
  assign _01533_ = lut_lookup_1_else_else_else_else_acc_itm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13448" *) { and_dcpl_403, and_dcpl_403, and_dcpl_403, and_dcpl_403, and_dcpl_403, and_dcpl_403, and_dcpl_403, and_dcpl_403, and_dcpl_403 };
  assign chn_lut_out_and_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5452" *) _02318_;
  assign and_dcpl_72 = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5453" *) main_stage_v_5;
  assign _01534_ = and_dcpl_72 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5453" *) lut_lookup_1_and_svs_2;
  assign chn_lut_out_and_13_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5454" *) _03352_;
  assign _01535_ = and_dcpl_72 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5455" *) lut_lookup_2_and_svs_2;
  assign chn_lut_out_and_14_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5456" *) _03353_;
  assign _01536_ = and_dcpl_72 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5457" *) lut_lookup_3_and_svs_2;
  assign chn_lut_out_and_15_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5458" *) _03354_;
  assign _01537_ = and_dcpl_72 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5459" *) lut_lookup_4_and_svs_2;
  assign chn_lut_out_and_16_cse = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5460" *) _03355_;
  assign lut_lookup_and_138_cse = _02319_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5461" *) lut_lookup_or_3_tmp;
  assign lut_lookup_and_139_cse = lut_lookup_unequal_tmp_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5462" *) lut_lookup_or_3_tmp;
  assign lut_lookup_and_136_cse = _02319_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5463" *) lut_lookup_or_7_tmp;
  assign lut_lookup_and_137_cse = lut_lookup_unequal_tmp_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5464" *) lut_lookup_or_7_tmp;
  assign lut_lookup_and_134_cse = _02319_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5465" *) lut_lookup_or_11_tmp;
  assign lut_lookup_and_135_cse = lut_lookup_unequal_tmp_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5466" *) lut_lookup_or_11_tmp;
  assign lut_lookup_and_132_cse = _02319_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5467" *) lut_lookup_or_15_tmp;
  assign lut_lookup_and_133_cse = lut_lookup_unequal_tmp_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5468" *) lut_lookup_or_15_tmp;
  assign cfg_precision_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5469" *) mux_580_cse;
  assign FpAdd_8U_23U_2_is_addition_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5471" *) _02320_;
  assign FpAdd_8U_23U_1_is_addition_and_1_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5472" *) _02100_;
  assign cfg_lut_le_index_offset_and_1_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5473" *) mux_tmp_10;
  assign _01538_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5483" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign and_284_rgt = _01538_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5483" *) _02321_;
  assign and_286_rgt = _01538_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5484" *) reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign and_288_rgt = and_524_rgt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5486" *) _02321_;
  assign and_290_rgt = and_524_rgt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5487" *) reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign FpAdd_8U_23U_2_and_35_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5488" *) _02322_;
  assign and_292_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5489" *) reg_lut_lookup_1_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign _01539_ = and_dcpl_540 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5495" *) reg_cfg_precision_1_sva_st_12_cse_1[1];
  assign and_961_cse = _01539_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5496" *) _02323_;
  assign IsNaN_8U_23U_3_aelse_and_3_cse = _00928_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5500" *) _02107_;
  assign and_300_rgt = _01538_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5501" *) _02324_;
  assign and_302_rgt = _01538_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5502" *) reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign and_304_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5503" *) _02325_;
  assign and_306_rgt = and_524_rgt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5504" *) reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign FpAdd_8U_23U_2_and_36_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5505" *) _02326_;
  assign and_308_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5506" *) reg_lut_lookup_2_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign and_316_rgt = _01538_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5510" *) _02327_;
  assign and_318_rgt = _01538_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5511" *) reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign and_320_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5512" *) _02328_;
  assign and_322_rgt = and_524_rgt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5513" *) reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign FpAdd_8U_23U_2_and_37_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5514" *) _02107_;
  assign and_324_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5515" *) reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign and_330_rgt = _01538_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5519" *) _02329_;
  assign and_332_rgt = _01538_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5520" *) reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign and_524_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5521" *) _02281_;
  assign and_334_rgt = and_524_rgt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5522" *) _02329_;
  assign and_336_rgt = and_524_rgt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5523" *) reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign and_338_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5524" *) reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign _00924_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5525" *) _02101_;
  assign cfg_lut_le_start_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5525" *) mux_tmp_35;
  assign _01540_ = nor_193_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5527" *) _02299_;
  assign and_344_rgt = _01540_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5527" *) or_cse;
  assign _01541_ = or_66_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5528" *) _02299_;
  assign and_347_rgt = _01541_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5529" *) or_cse;
  assign FpMantRNE_49U_24U_1_else_o_mant_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5538" *) mux_42_nl;
  assign and_355_m1c = or_dcpl_51 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5539" *) or_cse;
  assign FpAdd_8U_23U_o_expo_and_3_ssc = _02330_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5549" *) and_355_m1c;
  assign _01542_ = _02332_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5551" *) FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49];
  assign FpAdd_8U_23U_and_51_ssc = _01542_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5551" *) and_355_m1c;
  assign _01543_ = lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5553" *) FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49];
  assign FpAdd_8U_23U_and_43_ssc = _01543_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5553" *) and_355_m1c;
  assign _01544_ = nor_193_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5559" *) or_cse;
  assign IsNaN_8U_23U_3_aelse_and_6_cse = _01117_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5562" *) _02334_;
  assign FpMantRNE_49U_24U_1_else_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5563" *) _02334_;
  assign _01545_ = _02336_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5570" *) FpAdd_8U_23U_2_int_mant_p1_1_sva_3[49];
  assign FpAdd_8U_23U_2_and_4_rgt = _01545_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5570" *) _02101_;
  assign _01546_ = lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5572" *) FpAdd_8U_23U_2_int_mant_p1_1_sva_3[49];
  assign FpAdd_8U_23U_2_and_5_rgt = _01546_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5572" *) _02101_;
  assign _01547_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5575" *) FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse;
  assign FpAdd_8U_23U_2_is_inf_and_cse = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5575" *) mux_tmp_35;
  assign _01548_ = and_dcpl_98 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5577" *) _02299_;
  assign and_364_rgt = _01548_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5577" *) or_cse;
  assign FpMantRNE_49U_24U_1_else_o_mant_and_1_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5588" *) mux_92_nl;
  assign and_375_m1c = or_dcpl_57 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5589" *) or_cse;
  assign FpAdd_8U_23U_o_expo_and_2_ssc = _02337_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5599" *) and_375_m1c;
  assign _01549_ = _02339_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5601" *) FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49];
  assign FpAdd_8U_23U_and_53_ssc = _01549_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5601" *) and_375_m1c;
  assign _01550_ = lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5603" *) FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49];
  assign FpAdd_8U_23U_and_45_ssc = _01550_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5603" *) and_375_m1c;
  assign and_401_cse = and_dcpl_98 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5608" *) or_cse;
  assign _01551_ = _02341_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5615" *) FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49];
  assign FpAdd_8U_23U_2_and_10_rgt = _01551_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5615" *) _02101_;
  assign _01552_ = lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5617" *) FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49];
  assign FpAdd_8U_23U_2_and_11_rgt = _01552_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5617" *) _02101_;
  assign IsNaN_8U_23U_8_aelse_and_1_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5619" *) _02342_;
  assign FpMantRNE_49U_24U_1_else_o_mant_and_2_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5629" *) mux_141_nl;
  assign FpAdd_8U_23U_o_expo_and_1_ssc = _02344_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5639" *) and_375_m1c;
  assign _01553_ = _02346_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5641" *) FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49];
  assign FpAdd_8U_23U_and_55_ssc = _01553_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5641" *) and_375_m1c;
  assign _01554_ = lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5643" *) FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49];
  assign FpAdd_8U_23U_and_47_ssc = _01554_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5643" *) and_375_m1c;
  assign _01555_ = _02348_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5649" *) FpAdd_8U_23U_2_int_mant_p1_3_sva_3[49];
  assign FpAdd_8U_23U_2_and_16_rgt = _01555_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5649" *) _02101_;
  assign _01556_ = lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5651" *) FpAdd_8U_23U_2_int_mant_p1_3_sva_3[49];
  assign FpAdd_8U_23U_2_and_17_rgt = _01556_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5651" *) _02101_;
  assign FpMantRNE_49U_24U_1_else_o_mant_and_3_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5660" *) mux_177_nl;
  assign FpAdd_8U_23U_o_expo_and_ssc = _02349_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5670" *) and_375_m1c;
  assign _01557_ = _02351_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5672" *) FpAdd_8U_23U_1_int_mant_p1_sva_3[49];
  assign FpAdd_8U_23U_and_57_ssc = _01557_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5672" *) and_375_m1c;
  assign _01558_ = lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5674" *) FpAdd_8U_23U_1_int_mant_p1_sva_3[49];
  assign FpAdd_8U_23U_and_49_ssc = _01558_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5674" *) and_375_m1c;
  assign _01559_ = _02353_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5679" *) FpAdd_8U_23U_2_int_mant_p1_sva_3[49];
  assign FpAdd_8U_23U_2_and_22_rgt = _01559_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5679" *) _02101_;
  assign _01560_ = lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5681" *) FpAdd_8U_23U_2_int_mant_p1_sva_3[49];
  assign FpAdd_8U_23U_2_and_23_rgt = _01560_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5681" *) _02101_;
  assign and_428_rgt = and_896_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5682" *) or_cse;
  assign and_427_cse = or_1857_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5683" *) or_cse;
  assign and_tmp_83 = main_stage_v_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5688" *) or_tmp_314;
  assign lut_lookup_if_else_if_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5690" *) mux_220_nl;
  assign cfg_precision_and_24_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5691" *) mux_tmp_220;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5698" *) mux_222_nl;
  assign and_430_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5699" *) _02112_;
  assign _01561_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5700" *) cfg_lut_le_function_1_sva_st_41;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5705" *) _02356_;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_1_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5713" *) mux_234_nl;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_1_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5717" *) _02357_;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_2_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5726" *) mux_247_nl;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_2_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5729" *) _02358_;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_3_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5737" *) mux_259_nl;
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_3_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5740" *) _02359_;
  assign cfg_lut_hybrid_priority_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5741" *) mux_tmp_265;
  assign and_854_cse = or_1853_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5745" *) lut_lookup_else_if_lor_5_lpi_1_dfm_5;
  assign lut_lookup_else_if_oelse_1_and_1_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5747" *) _02360_;
  assign and_852_cse = cfg_lut_le_function_1_sva_st_42 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5748" *) main_stage_v_4;
  assign and_846_cse = lut_lookup_unequal_tmp_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5751" *) lut_lookup_if_1_lor_5_lpi_1_dfm_5;
  assign lut_lookup_if_1_oelse_1_and_4_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5754" *) _02361_;
  assign lut_lookup_if_1_oelse_1_and_5_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5756" *) _02362_;
  assign and_82_cse = lut_lookup_else_if_lor_6_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5760" *) or_492_cse;
  assign and_843_cse = cfg_lut_le_function_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5761" *) main_stage_v_5;
  assign and_839_cse = or_492_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5764" *) lut_lookup_else_if_lor_7_lpi_1_dfm_5;
  assign lut_lookup_else_if_oelse_1_and_4_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5768" *) _02363_;
  assign lut_lookup_if_1_oelse_1_and_8_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5772" *) _02364_;
  assign and_835_cse = or_492_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5775" *) lut_lookup_else_if_lor_1_lpi_1_dfm_5;
  assign _01562_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5776" *) _03449_;
  assign lut_lookup_le_uflow_and_cse = _01562_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5777" *) mux_tmp_265;
  assign lut_lookup_lo_index_0_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5782" *) mux_357_nl;
  assign and_465_cse = or_1202_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5783" *) and_dcpl_259;
  assign and_466_cse = nor_610_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5784" *) and_dcpl_259;
  assign lut_lookup_else_else_and_cse = _00918_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5791" *) mux_360_nl;
  assign and_832_cse = lut_lookup_unequal_tmp_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5792" *) main_stage_v_5;
  assign lut_lookup_lo_index_0_and_2_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5794" *) mux_366_nl;
  assign lut_lookup_lo_uflow_and_4_cse = _00961_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5797" *) mux_tmp_220;
  assign _01563_ = FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5799" *) or_cse;
  assign FpAdd_8U_23U_1_and_46_cse = _01102_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5801" *) _02366_;
  assign _01564_ = FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_1_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5803" *) or_cse;
  assign FpAdd_8U_23U_2_and_44_cse = _01109_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5805" *) _02100_;
  assign _01565_ = FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_2_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5807" *) or_cse;
  assign _01566_ = FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_3_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5809" *) or_cse;
  assign _01567_ = _02367_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5811" *) lut_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  assign _01568_ = and_dcpl_309 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5813" *) cfg_lut_le_function_rsci_d;
  assign _01569_ = _01568_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5813" *) or_cse;
  assign _01570_ = and_dcpl_309 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5814" *) _02368_;
  assign _01571_ = _01570_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5814" *) or_cse;
  assign _01572_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5814" *) _03453_;
  assign FpAdd_8U_23U_1_is_a_greater_oelse_and_cse = _01572_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5814" *) mux_580_cse;
  assign IsZero_8U_23U_4_and_cse = _01105_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5817" *) _02366_;
  assign _01573_ = _02369_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5819" *) lut_lookup_1_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  assign _01574_ = and_dcpl_309 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5821" *) or_cse;
  assign _01575_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5821" *) _03454_;
  assign FpAdd_8U_23U_2_is_a_greater_oelse_and_cse = _01575_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5821" *) mux_580_cse;
  assign _01576_ = _02370_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5823" *) lut_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  assign IsZero_8U_23U_4_and_1_cse = _01105_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5825" *) _02100_;
  assign _01577_ = _02371_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5827" *) lut_lookup_2_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  assign _01578_ = _02372_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5829" *) lut_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  assign _01579_ = _02373_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5831" *) lut_lookup_3_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  assign _01580_ = _02374_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5834" *) lut_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  assign _01581_ = _02375_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5836" *) lut_lookup_4_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  assign IsZero_8U_23U_7_and_3_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5837" *) _02103_;
  assign and_525_rgt = or_26_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5839" *) or_cse;
  assign _01582_ = and_956_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5841" *) or_cse;
  assign _01583_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5841" *) _03455_;
  assign IsNaN_8U_23U_1_aelse_and_4_cse = _01583_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5841" *) mux_tmp_10;
  assign _01584_ = and_956_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5843" *) _02281_;
  assign and_527_rgt = _01584_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5843" *) or_cse;
  assign _01585_ = and_956_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5844" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign and_529_rgt = _01585_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5844" *) or_cse;
  assign _01586_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5846" *) _03457_;
  assign IsNaN_8U_23U_1_aelse_and_5_cse = _01586_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5846" *) mux_tmp_10;
  assign and_551_rgt = mux_1185_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5851" *) or_cse;
  assign _01587_ = _02376_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5852" *) and_553_m1c;
  assign _01588_ = _02377_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5853" *) and_555_m1c;
  assign _01589_ = IsNaN_8U_23U_4_land_1_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5854" *) and_553_m1c;
  assign _01590_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5855" *) and_555_m1c;
  assign _01591_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5857" *) _02378_;
  assign _01592_ = _01591_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5857" *) reg_cfg_precision_1_sva_st_12_cse_1[1];
  assign and_562_m1c = _01592_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5857" *) and_dcpl_351;
  assign _01593_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5860" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
  assign _01594_ = _01593_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5861" *) reg_cfg_precision_1_sva_st_12_cse_1[1];
  assign and_559_rgt = _01594_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5861" *) and_dcpl_351;
  assign lut_lookup_and_126_rgt = _02379_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5862" *) and_562_m1c;
  assign lut_lookup_and_127_rgt = IsNaN_8U_23U_8_land_2_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5863" *) and_562_m1c;
  assign _01595_ = or_1688_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5865" *) main_stage_v_2;
  assign and_564_rgt = _01595_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5865" *) and_401_cse;
  assign and_567_m1c = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5867" *) _02380_;
  assign and_566_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5868" *) IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
  assign lut_lookup_and_124_rgt = _02381_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5869" *) and_567_m1c;
  assign lut_lookup_and_125_rgt = IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5870" *) and_567_m1c;
  assign _01596_ = and_dcpl_364 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5871" *) or_cse;
  assign and_572_m1c = _01596_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5871" *) _02380_;
  assign and_570_rgt = _01596_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5872" *) IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
  assign lut_lookup_and_122_rgt = _02379_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5873" *) and_572_m1c;
  assign lut_lookup_and_123_rgt = IsNaN_8U_23U_8_land_2_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5874" *) and_572_m1c;
  assign and_577_m1c = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5878" *) _02382_;
  assign and_576_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5879" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  assign lut_lookup_and_120_rgt = _02381_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5880" *) and_577_m1c;
  assign lut_lookup_and_121_rgt = IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5881" *) and_577_m1c;
  assign and_582_m1c = _01596_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5882" *) _02382_;
  assign and_580_rgt = _01596_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5883" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  assign lut_lookup_and_118_rgt = _02383_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5884" *) and_582_m1c;
  assign lut_lookup_and_119_rgt = nor_482_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5885" *) and_582_m1c;
  assign _01597_ = or_1688_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5887" *) and_dcpl_98;
  assign _01598_ = _01597_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5887" *) main_stage_v_2;
  assign and_586_rgt = _01598_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5887" *) or_cse;
  assign and_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5891" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign and_588_rgt = mux_1186_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5893" *) or_cse;
  assign _01599_ = _02384_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5894" *) and_590_m1c;
  assign _01600_ = _02385_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5895" *) and_592_m1c;
  assign _01601_ = IsNaN_8U_23U_4_land_lpi_1_dfm_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5896" *) and_590_m1c;
  assign _01602_ = IsNaN_8U_23U_1_land_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5897" *) and_592_m1c;
  assign and_597_m1c = _01596_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5898" *) _02386_;
  assign and_595_rgt = _01596_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5899" *) reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse;
  assign lut_lookup_and_112_rgt = _02387_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5900" *) and_597_m1c;
  assign lut_lookup_and_113_rgt = nor_469_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5901" *) and_597_m1c;
  assign _01603_ = and_896_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5902" *) cfg_lut_le_function_1_sva_st_41;
  assign and_604_rgt = _01603_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5902" *) or_cse;
  assign _01604_ = or_1857_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5903" *) _02112_;
  assign and_606_rgt = _01604_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5903" *) or_cse;
  assign lut_lookup_else_if_oelse_1_and_8_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5910" *) _02388_;
  assign and_826_cse = cfg_lut_le_function_1_sva_st_41 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5911" *) main_stage_v_3;
  assign and_120_nl = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5914" *) mux_tmp_704;
  assign lut_lookup_lo_index_0_and_4_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5916" *) mux_707_nl;
  assign lut_lookup_if_1_oelse_1_and_12_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5921" *) _02390_;
  assign lut_lookup_lo_index_0_and_6_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5923" *) mux_729_nl;
  assign lut_lookup_if_1_oelse_1_and_14_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5925" *) _02391_;
  assign lut_lookup_if_if_oelse_1_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5935" *) _02392_;
  assign mux_771_cse = mux_1281_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5943" *) _02112_;
  assign lut_lookup_if_else_if_and_4_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5949" *) mux_775_nl;
  assign lut_lookup_1_IntLog2_32U_and_nl = IntLog2_32U_ac_int_cctor_1_30_0_1_sva_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5955" *) lut_lookup_1_IntLog2_32U_acc_1_nl;
  assign and_649_nl = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5956" *) _02393_;
  assign and_1142_cse = _02058_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5962" *) _02033_;
  assign _01605_ = lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5982" *) or_tmp_314;
  assign _01606_ = _03905_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5989" *) or_cse;
  assign and_898_cse = _01606_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5990" *) core_wen;
  assign _01607_ = _02639_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5991" *) or_cse;
  assign and_901_cse = _01607_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5992" *) core_wen;
  assign and_905_cse = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5993" *) core_wen;
  assign and_814_cse = cfg_lut_le_function_1_sva_st_42 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5994" *) lut_lookup_else_unequal_tmp_18;
  assign _01608_ = FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5996" *) lut_lookup_else_else_slc_32_mdf_1_sva_7;
  assign and_132_nl = _01608_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5996" *) mux_tmp_704;
  assign mux_789_cse = mux_1280_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5998" *) cfg_lut_le_function_1_sva_st_41;
  assign and_134_cse = and_852_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5999" *) or_tmp_314;
  assign and_653_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6000" *) _02396_;
  assign and_1141_cse = _02060_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6010" *) _02034_;
  assign _01609_ = lut_lookup_2_if_else_slc_32_svs_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6014" *) mux_tmp_704;
  assign lut_lookup_2_IntLog2_32U_and_nl = IntLog2_32U_ac_int_cctor_1_30_0_2_sva_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6019" *) lut_lookup_2_IntLog2_32U_acc_1_nl;
  assign and_657_nl = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6020" *) _02398_;
  assign and_907_cse = and_905_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6025" *) or_1857_cse;
  assign _01610_ = lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6040" *) or_tmp_314;
  assign and_811_cse = cfg_lut_le_function_1_sva_st_42 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6046" *) lut_lookup_else_unequal_tmp_12;
  assign _01611_ = FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6048" *) lut_lookup_else_else_slc_32_mdf_2_sva_7;
  assign and_143_nl = _01611_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6048" *) mux_tmp_704;
  assign mux_845_cse = mux_1279_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6050" *) cfg_lut_le_function_1_sva_st_41;
  assign lut_lookup_else_else_and_5_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6054" *) mux_853_nl;
  assign and_661_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6055" *) _02400_;
  assign and_1140_cse = _02061_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6057" *) _02035_;
  assign _01612_ = lut_lookup_3_if_else_slc_32_svs_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6060" *) mux_tmp_704;
  assign lut_lookup_3_IntLog2_32U_and_nl = IntLog2_32U_ac_int_cctor_1_30_0_3_sva_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6065" *) lut_lookup_3_IntLog2_32U_acc_1_nl;
  assign and_665_nl = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6066" *) _02402_;
  assign _01613_ = FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6092" *) lut_lookup_else_else_slc_32_mdf_3_sva_7;
  assign and_153_nl = _01613_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6092" *) mux_tmp_704;
  assign mux_900_cse = mux_1278_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6094" *) cfg_lut_le_function_1_sva_st_41;
  assign and_668_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6095" *) _02404_;
  assign and_1139_cse = _02062_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6097" *) _02036_;
  assign lut_lookup_else_1_and_6_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6101" *) mux_919_nl;
  assign lut_lookup_4_IntLog2_32U_and_nl = IntLog2_32U_ac_int_cctor_1_30_0_sva_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6107" *) lut_lookup_4_IntLog2_32U_acc_1_nl;
  assign and_672_nl = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6108" *) _02405_;
  assign _01614_ = FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6133" *) lut_lookup_else_else_slc_32_mdf_sva_7;
  assign and_164_nl = _01614_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6133" *) mux_tmp_704;
  assign mux_959_cse = mux_1269_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6135" *) cfg_lut_le_function_1_sva_st_41;
  assign and_676_rgt = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6136" *) _02406_;
  assign and_1138_cse = _02063_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6138" *) _02037_;
  assign lut_lookup_else_and_8_cse = _00961_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6140" *) mux_tmp_978;
  assign and_679_rgt = nor_792_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6141" *) or_cse;
  assign and_42_cse = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6142" *) or_66_cse;
  assign and_178_cse = reg_cfg_lut_le_function_1_sva_st_20_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6144" *) mux_982_cse;
  assign and_1179_nl = mux_793_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6145" *) cfg_lut_le_function_1_sva_st_41;
  assign lut_lookup_else_else_and_9_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6147" *) mux_1004_nl;
  assign lut_lookup_else_1_and_9_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6149" *) mux_1053_nl;
  assign lut_lookup_lo_index_0_and_8_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6151" *) mux_1056_nl;
  assign and_795_cse = _02080_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6152" *) _02031_;
  assign and_794_cse = _02076_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6153" *) _02038_;
  assign and_789_cse = _02077_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6154" *) _02039_;
  assign and_787_cse = _02078_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6155" *) _02040_;
  assign and_784_cse = _02081_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6156" *) _02041_;
  assign IsNaN_8U_23U_8_and_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6162" *) mux_1067_nl;
  assign and_780_cse = _02079_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6163" *) _02032_;
  assign IsNaN_8U_23U_8_and_2_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6170" *) mux_1074_nl;
  assign lut_lookup_else_1_and_13_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6172" *) mux_1106_nl;
  assign lut_lookup_else_1_and_16_cse = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6174" *) mux_1115_nl;
  assign FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w0 = FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6210" *) _03528_;
  assign lut_lookup_1_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6216" *) _02042_;
  assign FpMantRNE_49U_24U_2_else_carry_1_sva_mx0w0 = FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6230" *) _03552_;
  assign lut_lookup_1_FpMantRNE_49U_24U_2_else_and_tmp = FpMantRNE_49U_24U_2_else_carry_1_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6232" *) _02043_;
  assign FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w0 = FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6250" *) _03576_;
  assign lut_lookup_2_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6256" *) _02044_;
  assign FpMantRNE_49U_24U_2_else_carry_2_sva_mx0w0 = FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6270" *) _03600_;
  assign lut_lookup_2_FpMantRNE_49U_24U_2_else_and_tmp = FpMantRNE_49U_24U_2_else_carry_2_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6272" *) _02045_;
  assign FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w0 = FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6290" *) _03624_;
  assign lut_lookup_3_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6296" *) _02046_;
  assign FpMantRNE_49U_24U_2_else_carry_3_sva_mx0w0 = FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6310" *) _03648_;
  assign lut_lookup_3_FpMantRNE_49U_24U_2_else_and_tmp = FpMantRNE_49U_24U_2_else_carry_3_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6312" *) _02047_;
  assign FpMantRNE_49U_24U_1_else_carry_sva_mx0w0 = FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6330" *) _03672_;
  assign lut_lookup_4_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6336" *) _02048_;
  assign FpMantRNE_49U_24U_2_else_carry_sva_mx0w0 = FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[24] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6350" *) _03696_;
  assign lut_lookup_4_FpMantRNE_49U_24U_2_else_and_tmp = FpMantRNE_49U_24U_2_else_carry_sva_mx0w0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6352" *) _02049_;
  assign IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp = _02070_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6475" *) _02051_;
  assign IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp = _02072_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6481" *) _02052_;
  assign FpAdd_8U_23U_and_59_nl = _02418_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6596" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c;
  assign _01615_ = FpAdd_8U_23U_1_and_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6598" *) _02419_;
  assign FpAdd_8U_23U_and_61_nl = _01615_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6598" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c;
  assign FpAdd_8U_23U_1_and_35_nl = FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6599" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c;
  assign FpAdd_8U_23U_and_35_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6600" *) _02393_;
  assign FpAdd_8U_23U_1_and_tmp = lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6607" *) reg_lut_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign FpAdd_8U_23U_2_and_nl = _02421_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6624" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_5_m1c;
  assign _01616_ = FpAdd_8U_23U_2_and_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6626" *) _02422_;
  assign FpAdd_8U_23U_2_and_6_nl = _01616_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6626" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_5_m1c;
  assign FpAdd_8U_23U_2_and_28_nl = FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6627" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_5_m1c;
  assign FpAdd_8U_23U_2_and_9_nl = IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6628" *) _02396_;
  assign FpAdd_8U_23U_2_and_tmp = lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6634" *) lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign FpAdd_8U_23U_and_63_nl = _02424_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6647" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c;
  assign _01617_ = FpAdd_8U_23U_1_and_1_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6649" *) _02425_;
  assign FpAdd_8U_23U_and_65_nl = _01617_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6649" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c;
  assign FpAdd_8U_23U_1_and_37_nl = FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6650" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c;
  assign FpAdd_8U_23U_and_37_nl = IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6651" *) _02398_;
  assign FpAdd_8U_23U_1_and_1_tmp = lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6658" *) reg_lut_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp = _02074_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6662" *) _02053_;
  assign FpAdd_8U_23U_2_and_29_nl = _02427_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6677" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_7_m1c;
  assign _01618_ = FpAdd_8U_23U_2_and_1_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6679" *) _02428_;
  assign FpAdd_8U_23U_2_and_13_nl = _01618_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6679" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_7_m1c;
  assign FpAdd_8U_23U_2_and_30_nl = FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6680" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_7_m1c;
  assign FpAdd_8U_23U_2_and_15_nl = IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6681" *) _02400_;
  assign FpAdd_8U_23U_2_and_1_tmp = lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6687" *) lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign FpAdd_8U_23U_and_67_nl = _02430_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6700" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c;
  assign _01619_ = FpAdd_8U_23U_1_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6702" *) _02431_;
  assign FpAdd_8U_23U_and_69_nl = _01619_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6702" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c;
  assign FpAdd_8U_23U_1_and_39_nl = FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6703" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c;
  assign FpAdd_8U_23U_and_39_nl = IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6704" *) _02402_;
  assign FpAdd_8U_23U_1_and_2_tmp = lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6711" *) reg_lut_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign FpAdd_8U_23U_2_and_31_nl = _02433_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6728" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_9_m1c;
  assign _01620_ = FpAdd_8U_23U_2_and_2_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6730" *) _02434_;
  assign FpAdd_8U_23U_2_and_19_nl = _01620_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6730" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_9_m1c;
  assign FpAdd_8U_23U_2_and_32_nl = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6731" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_9_m1c;
  assign FpAdd_8U_23U_2_and_21_nl = IsNaN_8U_23U_8_land_3_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6732" *) _02404_;
  assign FpAdd_8U_23U_2_and_2_tmp = lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6738" *) lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign FpAdd_8U_23U_and_71_nl = _02436_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6751" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c;
  assign _01621_ = FpAdd_8U_23U_1_and_3_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6753" *) _02437_;
  assign FpAdd_8U_23U_and_73_nl = _01621_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6753" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c;
  assign FpAdd_8U_23U_1_and_41_nl = FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6754" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c;
  assign FpAdd_8U_23U_and_41_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6755" *) _02405_;
  assign FpAdd_8U_23U_1_and_3_tmp = lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6762" *) reg_lut_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign FpAdd_8U_23U_2_and_33_nl = _02439_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6779" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_11_m1c;
  assign _01622_ = FpAdd_8U_23U_2_and_3_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6781" *) _02440_;
  assign FpAdd_8U_23U_2_and_25_nl = _01622_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6781" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_11_m1c;
  assign FpAdd_8U_23U_2_and_34_nl = FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6782" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_11_m1c;
  assign FpAdd_8U_23U_2_and_27_nl = IsNaN_8U_23U_8_land_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6783" *) _02406_;
  assign FpAdd_8U_23U_2_and_3_tmp = lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6789" *) lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse = lut_lookup_lo_miss_1_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6846" *) lut_lookup_le_miss_1_sva;
  assign lut_lookup_if_1_lut_lookup_if_1_and_11_nl = lut_lookup_if_1_else_lo_int_1_lpi_1_dfm_1[8] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6854" *) _00074_[34];
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_1_cse = lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6863" *) cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_cse = lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6865" *) cfg_lut_hybrid_priority_1_sva_10;
  assign _01623_ = lut_lookup_else_if_else_le_fra_1_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6871" *) { lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 };
  assign _01624_ = _01623_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6871" *) { _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34] };
  assign _01625_ = _01624_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6872" *) { lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3], lut_lookup_1_else_if_else_if_acc_nl[3] };
  assign lut_lookup_le_fraction_1_lpi_1_dfm_9 = _01625_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6872" *) { _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34] };
  assign _01626_ = lut_lookup_if_1_else_lo_int_1_lpi_1_dfm_1[7:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6889" *) { _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34] };
  assign lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_1 = _01626_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6890" *) { _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34] };
  assign _01627_ = lut_lookup_if_1_else_lo_fra_1_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6894" *) { lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 };
  assign _01628_ = _01627_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6894" *) { _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34] };
  assign _01629_ = _01628_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6895" *) { _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34] };
  assign lut_lookup_lo_fraction_1_lpi_1_dfm_1 = _01629_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6895" *) { _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34] };
  assign lut_lookup_1_else_2_and_svs = lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6897" *) lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse = lut_lookup_lo_miss_2_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6905" *) lut_lookup_le_miss_2_sva;
  assign lut_lookup_if_1_lut_lookup_if_1_and_12_nl = lut_lookup_if_1_else_lo_int_2_lpi_1_dfm_1[8] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6913" *) _00079_[34];
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_2_cse = lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6917" *) cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_3_cse = lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6921" *) cfg_lut_hybrid_priority_1_sva_10;
  assign _01630_ = lut_lookup_else_if_else_le_fra_2_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6929" *) { lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 };
  assign _01631_ = _01630_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6929" *) { _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34] };
  assign _01632_ = _01631_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6930" *) { lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3], lut_lookup_2_else_if_else_if_acc_nl[3] };
  assign lut_lookup_le_fraction_2_lpi_1_dfm_9 = _01632_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6930" *) { _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34] };
  assign _01633_ = lut_lookup_if_1_else_lo_int_2_lpi_1_dfm_1[7:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6947" *) { _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34] };
  assign lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_1 = _01633_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6948" *) { _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34] };
  assign _01634_ = lut_lookup_if_1_else_lo_fra_2_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6952" *) { lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 };
  assign _01635_ = _01634_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6952" *) { _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34] };
  assign _01636_ = _01635_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6953" *) { _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34] };
  assign lut_lookup_lo_fraction_2_lpi_1_dfm_1 = _01636_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6953" *) { _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34] };
  assign lut_lookup_2_else_2_and_svs = lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6955" *) lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse = lut_lookup_lo_miss_3_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6963" *) lut_lookup_le_miss_3_sva;
  assign lut_lookup_if_1_lut_lookup_if_1_and_13_nl = lut_lookup_if_1_else_lo_int_3_lpi_1_dfm_1[8] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6971" *) _00084_[34];
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_4_cse = lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6975" *) cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_5_cse = lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6979" *) cfg_lut_hybrid_priority_1_sva_10;
  assign _01637_ = lut_lookup_else_if_else_le_fra_3_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6987" *) { lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 };
  assign _01638_ = _01637_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6987" *) { _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34] };
  assign _01639_ = _01638_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6988" *) { lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3], lut_lookup_3_else_if_else_if_acc_nl[3] };
  assign lut_lookup_le_fraction_3_lpi_1_dfm_9 = _01639_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6988" *) { _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34] };
  assign _01640_ = lut_lookup_if_1_else_lo_int_3_lpi_1_dfm_1[7:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7005" *) { _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34] };
  assign lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_1 = _01640_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7006" *) { _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34] };
  assign _01641_ = lut_lookup_if_1_else_lo_fra_3_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7010" *) { lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 };
  assign _01642_ = _01641_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7010" *) { _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34] };
  assign _01643_ = _01642_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7011" *) { _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34] };
  assign lut_lookup_lo_fraction_3_lpi_1_dfm_1 = _01643_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7011" *) { _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34] };
  assign lut_lookup_3_else_2_and_svs = lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7013" *) lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0;
  assign lut_lookup_if_1_lut_lookup_if_1_and_14_nl = lut_lookup_if_1_else_lo_int_lpi_1_dfm_1[8] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7021" *) _00089_[34];
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_6_cse = lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7025" *) cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse = lut_lookup_lo_miss_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7027" *) lut_lookup_le_miss_sva;
  assign lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_7_cse = lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7037" *) cfg_lut_hybrid_priority_1_sva_10;
  assign _01644_ = lut_lookup_else_if_else_le_fra_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7045" *) { lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 };
  assign _01645_ = _01644_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7045" *) { _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34] };
  assign _01646_ = _01645_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7046" *) { lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3], lut_lookup_4_else_if_else_if_acc_nl[3] };
  assign lut_lookup_le_fraction_lpi_1_dfm_9 = _01646_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7046" *) { _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34] };
  assign _01647_ = lut_lookup_if_1_else_lo_int_lpi_1_dfm_1[7:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7063" *) { _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34] };
  assign lut_lookup_lo_index_0_7_0_lpi_1_dfm_1 = _01647_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7064" *) { _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34] };
  assign _01648_ = lut_lookup_if_1_else_lo_fra_sva_4 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7068" *) { lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2, lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 };
  assign _01649_ = _01648_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7068" *) { _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34] };
  assign _01650_ = _01649_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7069" *) { _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34] };
  assign lut_lookup_lo_fraction_lpi_1_dfm_1 = _01650_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7069" *) { _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34] };
  assign lut_lookup_4_else_2_and_svs = lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7071" *) lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0;
  assign _01651_ = reg_lut_lookup_if_unequal_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7075" *) _02208_;
  assign lut_lookup_and_5_cse = _01651_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7075" *) _02448_;
  assign _01652_ = _02319_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7077" *) cfg_lut_le_function_1_sva_10;
  assign lut_lookup_and_6_cse = _01652_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7077" *) _02448_;
  assign _01653_ = lut_lookup_unequal_tmp_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7079" *) cfg_lut_le_function_1_sva_10;
  assign lut_lookup_and_7_cse = _01653_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7079" *) _02448_;
  assign _01654_ = lut_lookup_le_miss_1_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7081" *) _02449_;
  assign _01655_ = cfg_lut_hybrid_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7083" *) _03730_;
  assign _01656_ = _03731_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7084" *) _02450_;
  assign _01657_ = cfg_lut_oflow_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7085" *) lut_lookup_1_else_2_and_svs;
  assign _01658_ = _01657_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7085" *) _02451_;
  assign _01659_ = cfg_lut_uflow_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7085" *) lut_lookup_1_and_svs_2;
  assign lut_lookup_and_13_cse = _01651_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7089" *) _02452_;
  assign _01660_ = _02453_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7091" *) cfg_lut_le_function_1_sva_10;
  assign lut_lookup_and_14_cse = _01660_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7091" *) _02452_;
  assign _01661_ = lut_lookup_else_unequal_tmp_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7093" *) cfg_lut_le_function_1_sva_10;
  assign lut_lookup_and_15_cse = _01661_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7093" *) _02452_;
  assign _01662_ = lut_lookup_le_miss_2_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7095" *) _02454_;
  assign _01663_ = cfg_lut_hybrid_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7097" *) _03734_;
  assign _01664_ = _03735_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7098" *) _02455_;
  assign _01665_ = cfg_lut_oflow_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7099" *) lut_lookup_2_else_2_and_svs;
  assign _01666_ = _01665_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7099" *) _02456_;
  assign _01667_ = cfg_lut_uflow_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7099" *) lut_lookup_2_and_svs_2;
  assign lut_lookup_and_21_cse = _01651_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7103" *) _02457_;
  assign lut_lookup_and_22_cse = _01660_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7105" *) _02457_;
  assign lut_lookup_and_23_cse = _01661_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7107" *) _02457_;
  assign _01668_ = lut_lookup_le_miss_3_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7109" *) _02458_;
  assign _01669_ = cfg_lut_hybrid_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7111" *) _03738_;
  assign _01670_ = _03739_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7112" *) _02459_;
  assign _01671_ = cfg_lut_oflow_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7113" *) lut_lookup_3_else_2_and_svs;
  assign _01672_ = _01671_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7113" *) _02460_;
  assign _01673_ = cfg_lut_uflow_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7113" *) lut_lookup_3_and_svs_2;
  assign lut_lookup_and_29_cse = _01651_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7117" *) _02461_;
  assign lut_lookup_and_30_cse = _01660_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7119" *) _02461_;
  assign lut_lookup_and_31_cse = _01661_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7121" *) _02461_;
  assign _01674_ = lut_lookup_le_miss_sva & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7123" *) _02462_;
  assign _01675_ = cfg_lut_hybrid_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7125" *) _03742_;
  assign _01676_ = _03743_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7126" *) _02463_;
  assign _01677_ = cfg_lut_oflow_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7127" *) lut_lookup_4_else_2_and_svs;
  assign _01678_ = _01677_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7127" *) _02464_;
  assign _01679_ = cfg_lut_uflow_priority_1_sva_10 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7127" *) lut_lookup_4_and_svs_2;
  assign main_stage_en_1 = chn_lut_in_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7128" *) or_cse;
  assign FpNormalize_8U_49U_oelse_not_9 = _02082_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7380" *) lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl[8];
  assign FpNormalize_8U_49U_2_oelse_not_9 = _02083_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7386" *) lut_lookup_1_FpNormalize_8U_49U_2_acc_nl[8];
  assign FpNormalize_8U_49U_oelse_not_11 = _02084_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7392" *) lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl[8];
  assign FpNormalize_8U_49U_2_oelse_not_11 = _02085_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7398" *) lut_lookup_2_FpNormalize_8U_49U_2_acc_nl[8];
  assign FpNormalize_8U_49U_oelse_not_13 = _02086_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7404" *) lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl[8];
  assign FpNormalize_8U_49U_2_oelse_not_13 = _02087_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7410" *) lut_lookup_3_FpNormalize_8U_49U_2_acc_nl[8];
  assign FpNormalize_8U_49U_oelse_not_15 = _02088_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7416" *) lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl[8];
  assign FpNormalize_8U_49U_2_oelse_not_15 = _02089_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7422" *) lut_lookup_4_FpNormalize_8U_49U_2_acc_nl[8];
  assign _01680_ = reg_cfg_precision_1_sva_st_12_cse_1[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7468" *) main_stage_v_1;
  assign _01681_ = reg_cfg_precision_1_sva_st_13_cse_1[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7478" *) main_stage_v_2;
  assign _01682_ = FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7482" *) main_stage_v_3;
  assign and_tmp_5 = _01682_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7482" *) or_1857_cse;
  assign and_tmp_6 = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7483" *) or_1857_cse;
  assign _01683_ = IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7487" *) lut_lookup_else_1_slc_32_mdf_1_sva_6;
  assign nor_tmp_12 = _01683_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7487" *) main_stage_v_2;
  assign nor_tmp_14 = lut_lookup_else_1_slc_32_mdf_1_sva_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7488" *) FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5;
  assign _01684_ = IsNaN_8U_23U_8_land_1_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7490" *) main_stage_v_2;
  assign _01685_ = IsNaN_8U_23U_8_land_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7498" *) main_stage_v_3;
  assign nor_tmp_32 = _01257_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7506" *) main_stage_v_2;
  assign nor_tmp_34 = lut_lookup_else_1_slc_32_mdf_2_sva_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7507" *) FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5;
  assign _01686_ = lut_lookup_2_FpMantRNE_49U_24U_2_else_and_tmp & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7509" *) main_stage_v_2;
  assign _01687_ = _01686_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7509" *) and_dcpl_98;
  assign _01688_ = FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7515" *) main_stage_v_3;
  assign and_tmp_14 = _01688_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7515" *) or_1857_cse;
  assign _01689_ = IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7517" *) lut_lookup_else_1_slc_32_mdf_3_sva_6;
  assign nor_tmp_44 = _01689_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7517" *) main_stage_v_2;
  assign _01690_ = FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7519" *) main_stage_v_3;
  assign and_tmp_19 = _01690_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7519" *) or_1857_cse;
  assign nor_tmp_57 = lut_lookup_else_1_slc_32_mdf_sva_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7522" *) FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5;
  assign _01691_ = lut_lookup_1_if_else_slc_32_svs_st_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7528" *) main_stage_v_4;
  assign _01692_ = _01691_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7529" *) or_tmp_314;
  assign _01693_ = FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7533" *) main_stage_v_3;
  assign and_tmp_27 = _01693_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7533" *) or_1857_cse;
  assign _01694_ = lut_lookup_2_if_else_slc_32_svs_st_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7534" *) main_stage_v_4;
  assign _01695_ = _01694_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7535" *) or_tmp_314;
  assign _01696_ = lut_lookup_3_if_else_slc_32_svs_st_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7538" *) main_stage_v_4;
  assign _01697_ = _01696_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7539" *) or_tmp_314;
  assign _01698_ = and_852_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7541" *) _02054_;
  assign _01699_ = lut_lookup_4_if_else_slc_32_svs_st_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7545" *) main_stage_v_4;
  assign _01700_ = _01699_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7546" *) or_tmp_314;
  assign _01701_ = _03769_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7552" *) lut_lookup_else_if_lor_5_lpi_1_dfm_6;
  assign _01702_ = cfg_precision_1_sva_st_72[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7561" *) cfg_lut_le_function_1_sva_10;
  assign _01703_ = _01702_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7561" *) main_stage_v_5;
  assign _01704_ = lut_lookup_unequal_tmp_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7565" *) lut_lookup_if_1_lor_6_lpi_1_dfm_5;
  assign _01705_ = or_1851_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7571" *) lut_lookup_else_if_lor_7_lpi_1_dfm_6;
  assign and_850_cse = lut_lookup_unequal_tmp_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7573" *) lut_lookup_if_1_lor_7_lpi_1_dfm_5;
  assign _01706_ = or_1851_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7576" *) lut_lookup_else_if_lor_1_lpi_1_dfm_6;
  assign and_848_cse = lut_lookup_unequal_tmp_13 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7578" *) lut_lookup_if_1_lor_1_lpi_1_dfm_5;
  assign nor_tmp_112 = lut_lookup_else_unequal_tmp_18 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7582" *) main_stage_v_4;
  assign and_dcpl_364 = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7588" *) and_956_cse;
  assign _01707_ = FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7604" *) or_cse;
  assign _01708_ = and_868_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7611" *) main_stage_v_2;
  assign and_tmp_59 = _01708_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7611" *) or_66_cse;
  assign _01709_ = IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7612" *) or_66_cse;
  assign and_tmp_61 = _01709_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7612" *) main_stage_v_2;
  assign _01710_ = IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7615" *) main_stage_v_2;
  assign and_tmp_69 = _01710_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7615" *) or_66_cse;
  assign _01711_ = lut_lookup_else_else_else_asn_mdf_1_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7625" *) cfg_lut_le_function_1_sva_st_41;
  assign _01712_ = _01711_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7625" *) FpAdd_8U_23U_1_mux_13_itm_4;
  assign _01713_ = _01712_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7625" *) lut_lookup_else_else_slc_32_mdf_1_sva_7;
  assign _01714_ = _01713_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7626" *) FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6;
  assign _01715_ = _01714_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7626" *) main_stage_v_3;
  assign and_tmp_92 = _01715_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7626" *) or_1857_cse;
  assign _01716_ = cfg_lut_le_function_1_sva_st_42 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7628" *) IsNaN_8U_23U_6_land_1_lpi_1_dfm_6;
  assign _01717_ = _01716_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7628" *) lut_lookup_else_else_slc_32_mdf_1_sva_8;
  assign nor_tmp_238 = _01717_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7628" *) main_stage_v_4;
  assign _01718_ = nor_tmp_14 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7631" *) main_stage_v_3;
  assign and_tmp_97 = _01718_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7631" *) or_1857_cse;
  assign _01719_ = lut_lookup_else_1_slc_32_mdf_1_sva_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7635" *) IsNaN_8U_23U_10_land_1_lpi_1_dfm_5;
  assign _01720_ = _01719_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7635" *) main_stage_v_4;
  assign and_tmp_98 = _01720_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7635" *) or_tmp_314;
  assign _01721_ = lut_lookup_else_else_else_asn_mdf_2_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7637" *) cfg_lut_le_function_1_sva_st_41;
  assign _01722_ = _01721_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7637" *) FpAdd_8U_23U_1_mux_29_itm_4;
  assign _01723_ = _01722_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7637" *) FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6;
  assign _01724_ = _01723_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7638" *) lut_lookup_else_else_slc_32_mdf_2_sva_7;
  assign _01725_ = _01724_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7638" *) main_stage_v_3;
  assign and_tmp_103 = _01725_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7638" *) or_1857_cse;
  assign _01726_ = cfg_lut_le_function_1_sva_st_42 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7640" *) IsNaN_8U_23U_6_land_2_lpi_1_dfm_6;
  assign _01727_ = _01726_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7640" *) lut_lookup_else_else_slc_32_mdf_2_sva_8;
  assign nor_tmp_260 = _01727_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7640" *) main_stage_v_4;
  assign _01728_ = lut_lookup_else_1_slc_32_mdf_2_sva_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *) main_stage_v_3;
  assign _01729_ = FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *) _02487_;
  assign _01730_ = lut_lookup_else_1_slc_32_mdf_2_sva_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7644" *) IsNaN_8U_23U_10_land_2_lpi_1_dfm_5;
  assign _01731_ = _01730_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7644" *) main_stage_v_4;
  assign and_tmp_108 = _01731_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7644" *) or_tmp_314;
  assign _01732_ = lut_lookup_else_else_else_asn_mdf_3_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7646" *) cfg_lut_le_function_1_sva_st_41;
  assign _01733_ = _01732_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7646" *) FpAdd_8U_23U_1_mux_45_itm_4;
  assign _01734_ = _01733_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7646" *) lut_lookup_else_else_slc_32_mdf_3_sva_7;
  assign _01735_ = _01734_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7647" *) FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6;
  assign _01736_ = _01735_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7647" *) main_stage_v_3;
  assign and_tmp_113 = _01736_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7647" *) or_1857_cse;
  assign _01737_ = cfg_lut_le_function_1_sva_st_42 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7649" *) IsNaN_8U_23U_6_land_3_lpi_1_dfm_6;
  assign _01738_ = _01737_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7649" *) lut_lookup_else_else_slc_32_mdf_3_sva_8;
  assign nor_tmp_281 = _01738_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7649" *) main_stage_v_4;
  assign _01739_ = lut_lookup_else_1_slc_32_mdf_3_sva_7 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7652" *) and_tmp_6;
  assign _01740_ = lut_lookup_else_1_slc_32_mdf_3_sva_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7654" *) IsNaN_8U_23U_10_land_3_lpi_1_dfm_5;
  assign _01741_ = _01740_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7654" *) main_stage_v_4;
  assign and_tmp_119 = _01741_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7654" *) or_tmp_314;
  assign _01742_ = lut_lookup_else_else_else_asn_mdf_sva_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7656" *) cfg_lut_le_function_1_sva_st_41;
  assign _01743_ = _01742_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7656" *) FpAdd_8U_23U_1_mux_61_itm_4;
  assign _01744_ = _01743_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7656" *) FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6;
  assign _01745_ = _01744_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7657" *) lut_lookup_else_else_slc_32_mdf_sva_7;
  assign _01746_ = _01745_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7657" *) main_stage_v_3;
  assign and_tmp_124 = _01746_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7657" *) or_1857_cse;
  assign and_tmp_130 = nor_tmp_57 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7659" *) and_tmp_6;
  assign _01747_ = lut_lookup_else_1_slc_32_mdf_sva_8 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7663" *) IsNaN_8U_23U_10_land_lpi_1_dfm_5;
  assign _01748_ = _01747_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7663" *) main_stage_v_4;
  assign and_tmp_131 = _01748_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7663" *) or_tmp_314;
  assign _01749_ = _01232_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7667" *) main_stage_v_2;
  assign _01750_ = _01749_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7667" *) or_66_cse;
  assign mux_tmp_1104 = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7671" *) or_26_cse;
  assign and_tmp_178 = chn_lut_in_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7673" *) or_1495_cse;
  assign and_dcpl_54 = _02490_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7674" *) reg_chn_lut_out_rsci_ld_core_psct_cse;
  assign and_dcpl_59 = and_dcpl_72 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7675" *) _02451_;
  assign and_dcpl_63 = and_dcpl_72 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7676" *) _02456_;
  assign and_dcpl_67 = and_dcpl_72 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7677" *) _02460_;
  assign and_dcpl_71 = and_dcpl_72 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7678" *) _02464_;
  assign _01751_ = _00010_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7680" *) chn_lut_out_rsci_bawt;
  assign and_dcpl_74 = _01751_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7680" *) reg_chn_lut_out_rsci_ld_core_psct_cse;
  assign and_dcpl_148 = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7684" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign and_dcpl_161 = or_66_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7686" *) or_cse;
  assign and_dcpl_162 = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7687" *) _02299_;
  assign and_dcpl_258 = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7720" *) cfg_lut_le_function_1_sva_st_42;
  assign and_dcpl_259 = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7721" *) _02201_;
  assign _01752_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7722" *) _02499_;
  assign and_dcpl_280 = _01752_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7723" *) _03815_;
  assign _01753_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7725" *) _03816_;
  assign and_dcpl_284 = _01753_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7725" *) _02502_;
  assign _01754_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7727" *) _03817_;
  assign and_dcpl_288 = _01754_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7727" *) _02504_;
  assign _01755_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7729" *) _03818_;
  assign and_dcpl_292 = _01755_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7729" *) _02506_;
  assign _01756_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7731" *) _03819_;
  assign and_dcpl_296 = _01756_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7731" *) _02508_;
  assign _01757_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7733" *) _03820_;
  assign and_dcpl_300 = _01757_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7733" *) _02510_;
  assign _01758_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7734" *) _02511_;
  assign and_dcpl_304 = _01758_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7735" *) _03821_;
  assign _01759_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7737" *) _03822_;
  assign and_dcpl_308 = _01759_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7737" *) _02514_;
  assign and_dcpl_314 = or_1495_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7739" *) or_cse;
  assign and_dcpl_315 = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7740" *) cfg_lut_le_function_rsci_d;
  assign and_dcpl_316 = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7741" *) _02368_;
  assign and_dcpl_351 = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7742" *) _02515_;
  assign _01760_ = or_1857_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7744" *) cfg_lut_le_function_1_sva_st_41;
  assign and_dcpl_403 = _01760_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7744" *) or_cse;
  assign _01761_ = and_896_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7745" *) _02112_;
  assign and_dcpl_405 = _01761_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7745" *) or_cse;
  assign or_tmp_1628 = main_stage_en_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7746" *) fsm_output[1];
  assign _01762_ = main_stage_v_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7748" *) _02280_;
  assign main_stage_v_1_mx0c1 = _01762_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7748" *) or_cse;
  assign _01763_ = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7749" *) _00033_;
  assign main_stage_v_2_mx0c1 = _01763_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7749" *) or_cse;
  assign _01764_ = main_stage_v_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7750" *) _00000_;
  assign main_stage_v_3_mx0c1 = _01764_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7750" *) or_cse;
  assign _01765_ = _00001_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7751" *) main_stage_v_4;
  assign main_stage_v_4_mx0c1 = _01765_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7751" *) or_cse;
  assign _01766_ = main_stage_v_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7752" *) _00032_;
  assign main_stage_v_5_mx0c1 = _01766_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7752" *) or_cse;
  assign _01767_ = lut_lookup_lo_uflow_1_lpi_1_dfm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7754" *) mux_tmp_1130;
  assign lut_lookup_else_2_else_else_if_mux_5_itm_1_mx0c1 = mux_1141_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7757" *) or_cse;
  assign _01768_ = lut_lookup_lo_uflow_2_lpi_1_dfm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7759" *) mux_tmp_1143;
  assign lut_lookup_else_2_else_else_if_mux_12_itm_1_mx0c1 = mux_1154_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7762" *) or_cse;
  assign _01769_ = lut_lookup_lo_uflow_3_lpi_1_dfm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7764" *) mux_tmp_1156;
  assign lut_lookup_else_2_else_else_if_mux_19_itm_1_mx0c1 = mux_1167_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7767" *) or_cse;
  assign _01770_ = lut_lookup_lo_uflow_lpi_1_dfm_3 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7769" *) mux_tmp_1169;
  assign lut_lookup_else_2_else_else_if_mux_26_itm_1_mx0c1 = mux_1180_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7772" *) or_cse;
  assign _01771_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7813" *) _02377_;
  assign and_553_m1c = _01771_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7813" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign and_555_m1c = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7814" *) _02528_;
  assign _01772_ = reg_cfg_lut_le_function_1_sva_st_19_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7816" *) _02385_;
  assign and_590_m1c = _01772_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7816" *) or_cse;
  assign and_592_m1c = _02529_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7818" *) or_cse;
  assign chn_lut_out_rsci_oswt_unreg = chn_lut_out_rsci_bawt & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7820" *) reg_chn_lut_out_rsci_ld_core_psct_cse;
  assign and_dcpl_540 = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7821" *) main_stage_v_1;
  assign and_dcpl_576 = main_stage_v_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7824" *) core_wen;
  assign and_dcpl_648 = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7845" *) main_stage_v_3;
  assign and_tmp_201 = lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7871" *) mux_tmp_1257;
  assign FpAdd_8U_23U_b_right_shift_qif_and_tmp = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7872" *) FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_cse;
  assign FpAdd_8U_23U_2_b_right_shift_qif_and_tmp = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7873" *) FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_3_cse;
  assign FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_1 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7874" *) FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_cse;
  assign FpAdd_8U_23U_b_right_shift_qif_and_tmp_1 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7875" *) FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_3_cse;
  assign FpAdd_8U_23U_b_right_shift_qif_and_tmp_2 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7876" *) FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_1_cse;
  assign FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_2 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7877" *) FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_2_cse;
  assign FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_3 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7878" *) FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_1_cse;
  assign FpAdd_8U_23U_b_right_shift_qif_and_tmp_3 = fsm_output[1] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7879" *) FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_2_cse;
  assign _01773_ = _02483_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7886" *) fsm_output[1];
  assign _01774_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7894" *) chn_lut_in_rsci_ld_core_psct_mx0c0;
  assign _01775_ = lut_lookup_else_2_mux_1_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7960" *) _02451_;
  assign _01776_ = lut_lookup_else_2_mux_27_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7961" *) _02456_;
  assign _01777_ = lut_lookup_else_2_mux_53_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7962" *) _02460_;
  assign _01778_ = lut_lookup_else_2_mux_79_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7963" *) _02464_;
  assign _01779_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8086" *) _03852_;
  assign _01780_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8094" *) _03853_;
  assign _01781_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8139" *) _02366_;
  assign _01782_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8224" *) main_stage_v_1;
  assign _01783_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8224" *) _03857_;
  assign _01784_ = and_dcpl_540 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8268" *) _02515_;
  assign _01785_ = _01784_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8269" *) or_cse;
  assign _01786_ = _01785_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8269" *) reg_cfg_precision_1_sva_st_12_cse_1[1];
  assign _01787_ = FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8278" *) _02281_;
  assign _01788_ = _03858_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8278" *) and_dcpl_540;
  assign _01789_ = _01788_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8278" *) or_cse;
  assign _01790_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8287" *) _03861_;
  assign _01791_ = _01790_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8287" *) not_tmp_47;
  assign _01792_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8310" *) _02552_;
  assign _01793_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8311" *) _03862_;
  assign _01794_ = _01793_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8311" *) _02322_;
  assign _01795_ = FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8333" *) _02281_;
  assign _01796_ = _03863_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8333" *) and_dcpl_540;
  assign _01797_ = _01796_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8333" *) or_cse;
  assign _01798_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8342" *) _03866_;
  assign _01799_ = _01798_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8342" *) _02107_;
  assign _01800_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8363" *) _02553_;
  assign _01801_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8364" *) _03867_;
  assign _01802_ = _01801_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8364" *) _02326_;
  assign _01803_ = _02281_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8373" *) FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5;
  assign _01804_ = _03868_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8374" *) and_dcpl_540;
  assign _01805_ = _01804_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8374" *) or_cse;
  assign _01806_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8383" *) _03871_;
  assign _01807_ = _01806_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8383" *) _02107_;
  assign _01808_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8412" *) _02554_;
  assign _01809_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8413" *) _03872_;
  assign _01810_ = _01809_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8413" *) _02107_;
  assign _01811_ = _02281_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8422" *) FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5;
  assign _01812_ = _03873_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8423" *) and_dcpl_540;
  assign _01813_ = _01812_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8423" *) or_cse;
  assign _01814_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8432" *) _03876_;
  assign _01815_ = _01814_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8432" *) _02107_;
  assign _01816_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8443" *) _02555_;
  assign _01817_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8444" *) _03877_;
  assign _01818_ = _01817_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8444" *) _02107_;
  assign _01819_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8453" *) main_stage_v_2;
  assign _01820_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8453" *) _03878_;
  assign _01821_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8503" *) _03880_;
  assign _01822_ = _01821_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8504" *) _02557_;
  assign _01823_ = _02558_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8515" *) core_wen;
  assign _01824_ = or_66_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8525" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign _01825_ = _01824_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8525" *) or_cse;
  assign _01826_ = _01825_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8526" *) _02559_;
  assign _01827_ = _01826_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8526" *) and_dcpl_576;
  assign _01828_ = or_1936_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8547" *) and_dcpl_576;
  assign _01829_ = _01828_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8548" *) reg_cfg_precision_1_sva_st_13_cse_1[1];
  assign _01830_ = _01829_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8548" *) nor_865_cse;
  assign _01831_ = _02560_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8558" *) and_dcpl_576;
  assign _01832_ = _01831_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8558" *) or_cse;
  assign _01833_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8568" *) FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_6_cse;
  assign _01834_ = _01833_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8568" *) mux_59_nl;
  assign _01835_ = _01833_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8645" *) mux_tmp_35;
  assign _01836_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8655" *) mux_61_nl;
  assign _01837_ = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8665" *) mux_66_nl;
  assign _01838_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8676" *) _03883_;
  assign _01839_ = _01838_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8676" *) _02561_;
  assign _01840_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8687" *) _02562_;
  assign _01841_ = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8696" *) mux_86_nl;
  assign _01842_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8723" *) IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_8_cse;
  assign _01843_ = _01842_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8724" *) _02563_;
  assign _01844_ = _02564_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8735" *) core_wen;
  assign _01845_ = or_66_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8745" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _01846_ = _01845_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8745" *) or_cse;
  assign _01847_ = _01846_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8746" *) _02565_;
  assign _01848_ = _01847_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8746" *) and_dcpl_576;
  assign _01849_ = _02673_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8768" *) and_dcpl_576;
  assign _01850_ = _01849_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8768" *) reg_cfg_precision_1_sva_st_13_cse_1[1];
  assign _01851_ = _01850_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8768" *) nor_865_cse;
  assign _01852_ = _02566_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8778" *) and_dcpl_576;
  assign _01853_ = _01852_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8778" *) or_cse;
  assign _01854_ = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8788" *) mux_121_nl;
  assign _01855_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8814" *) mux_123_nl;
  assign _01856_ = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8824" *) mux_128_nl;
  assign _01857_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8835" *) _03886_;
  assign _01858_ = _01857_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8836" *) _02567_;
  assign _01859_ = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8862" *) mux_135_nl;
  assign _01860_ = _01842_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8872" *) _02568_;
  assign _01861_ = _02569_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8883" *) core_wen;
  assign _01862_ = or_66_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8893" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign _01863_ = _01862_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8893" *) or_cse;
  assign _01864_ = _01863_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8894" *) _02570_;
  assign _01865_ = _01864_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8894" *) and_dcpl_576;
  assign _01866_ = _03890_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8916" *) and_dcpl_576;
  assign _01867_ = _01866_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8917" *) reg_cfg_precision_1_sva_st_13_cse_1[1];
  assign _01868_ = _01867_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8917" *) nor_865_cse;
  assign _01869_ = _02572_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8927" *) and_dcpl_576;
  assign _01870_ = _01869_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8927" *) or_cse;
  assign _01871_ = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8937" *) mux_157_nl;
  assign _01872_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8948" *) mux_159_nl;
  assign _01873_ = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8958" *) mux_164_nl;
  assign _01874_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8969" *) _03892_;
  assign _01875_ = _01874_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8970" *) _02573_;
  assign _01876_ = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8982" *) mux_171_nl;
  assign _01877_ = _01842_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8992" *) _02574_;
  assign _01878_ = _02575_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9003" *) core_wen;
  assign _01879_ = or_66_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9013" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _01880_ = _01879_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9013" *) or_cse;
  assign _01881_ = _01880_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9014" *) _02576_;
  assign _01882_ = _01881_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9014" *) and_dcpl_576;
  assign _01883_ = _03896_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9036" *) and_dcpl_576;
  assign _01884_ = _01883_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9037" *) reg_cfg_precision_1_sva_st_13_cse_1[1];
  assign _01885_ = _01884_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9037" *) nor_865_cse;
  assign _01886_ = _02578_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9047" *) and_dcpl_576;
  assign _01887_ = _01886_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9047" *) or_cse;
  assign _01888_ = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9057" *) mux_200_nl;
  assign _01889_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9068" *) mux_202_nl;
  assign _01890_ = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9078" *) mux_207_nl;
  assign _01891_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9089" *) _03898_;
  assign _01892_ = _01891_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9090" *) _02579_;
  assign _01893_ = _01547_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9102" *) mux_215_nl;
  assign _01894_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9111" *) main_stage_v_3;
  assign _01895_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9111" *) _03899_;
  assign _00961_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9129" *) lut_lookup_if_else_else_else_else_if_lut_lookup_if_else_else_else_else_if_or_3_cse;
  assign _01896_ = _00961_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9129" *) _02581_;
  assign _01897_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9139" *) mux_219_nl;
  assign _01898_ = lut_lookup_4_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9185" *) { lut_lookup_4_if_else_else_else_if_acc_nl[3], lut_lookup_4_if_else_else_else_if_acc_nl[3], lut_lookup_4_if_else_else_else_if_acc_nl[3], lut_lookup_4_if_else_else_else_if_acc_nl[3], lut_lookup_4_if_else_else_else_if_acc_nl[3], lut_lookup_4_if_else_else_else_if_acc_nl[3] };
  assign _01899_ = _01898_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9185" *) { _02582_, _02582_, _02582_, _02582_, _02582_, _02582_ };
  assign _01900_ = _01899_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9186" *) { lut_lookup_4_if_else_slc_32_svs_7, lut_lookup_4_if_else_slc_32_svs_7, lut_lookup_4_if_else_slc_32_svs_7, lut_lookup_4_if_else_slc_32_svs_7, lut_lookup_4_if_else_slc_32_svs_7, lut_lookup_4_if_else_slc_32_svs_7 };
  assign _01901_ = lut_lookup_3_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9191" *) { lut_lookup_3_if_else_else_else_if_acc_nl[3], lut_lookup_3_if_else_else_else_if_acc_nl[3], lut_lookup_3_if_else_else_else_if_acc_nl[3], lut_lookup_3_if_else_else_else_if_acc_nl[3], lut_lookup_3_if_else_else_else_if_acc_nl[3], lut_lookup_3_if_else_else_else_if_acc_nl[3] };
  assign _01902_ = _01901_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9191" *) { _02583_, _02583_, _02583_, _02583_, _02583_, _02583_ };
  assign _01903_ = _01902_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9192" *) { lut_lookup_3_if_else_slc_32_svs_7, lut_lookup_3_if_else_slc_32_svs_7, lut_lookup_3_if_else_slc_32_svs_7, lut_lookup_3_if_else_slc_32_svs_7, lut_lookup_3_if_else_slc_32_svs_7, lut_lookup_3_if_else_slc_32_svs_7 };
  assign _01904_ = lut_lookup_2_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9197" *) { lut_lookup_2_if_else_else_else_if_acc_nl[3], lut_lookup_2_if_else_else_else_if_acc_nl[3], lut_lookup_2_if_else_else_else_if_acc_nl[3], lut_lookup_2_if_else_else_else_if_acc_nl[3], lut_lookup_2_if_else_else_else_if_acc_nl[3], lut_lookup_2_if_else_else_else_if_acc_nl[3] };
  assign _01905_ = _01904_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9197" *) { _02584_, _02584_, _02584_, _02584_, _02584_, _02584_ };
  assign _01906_ = _01905_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9198" *) { lut_lookup_2_if_else_slc_32_svs_7, lut_lookup_2_if_else_slc_32_svs_7, lut_lookup_2_if_else_slc_32_svs_7, lut_lookup_2_if_else_slc_32_svs_7, lut_lookup_2_if_else_slc_32_svs_7, lut_lookup_2_if_else_slc_32_svs_7 };
  assign _01907_ = lut_lookup_1_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9203" *) { lut_lookup_1_if_else_else_else_if_acc_nl[3], lut_lookup_1_if_else_else_else_if_acc_nl[3], lut_lookup_1_if_else_else_else_if_acc_nl[3], lut_lookup_1_if_else_else_else_if_acc_nl[3], lut_lookup_1_if_else_else_else_if_acc_nl[3], lut_lookup_1_if_else_else_else_if_acc_nl[3] };
  assign _01908_ = _01907_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9203" *) { _02113_, _02113_, _02113_, _02113_, _02113_, _02113_ };
  assign _01909_ = _01908_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9204" *) { lut_lookup_1_if_else_slc_32_svs_7, lut_lookup_1_if_else_slc_32_svs_7, lut_lookup_1_if_else_slc_32_svs_7, lut_lookup_1_if_else_slc_32_svs_7, lut_lookup_1_if_else_slc_32_svs_7, lut_lookup_1_if_else_slc_32_svs_7 };
  assign _01910_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9223" *) FpAdd_8U_23U_1_lut_lookup_else_else_else_or_3_cse;
  assign _01911_ = _01910_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9224" *) mux_225_nl;
  assign _01912_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9244" *) mux_228_nl;
  assign _01913_ = _00961_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9255" *) _02587_;
  assign _01914_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9265" *) mux_232_nl;
  assign _01915_ = _01910_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9284" *) mux_237_nl;
  assign _01916_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9304" *) mux_240_nl;
  assign _01917_ = _00961_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9315" *) _02588_;
  assign _01918_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9325" *) mux_245_nl;
  assign _01919_ = _01910_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9344" *) mux_250_nl;
  assign _01920_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9364" *) mux_253_nl;
  assign _01921_ = _00961_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9375" *) _02589_;
  assign _01922_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9385" *) mux_257_nl;
  assign _01923_ = _01910_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9404" *) mux_262_nl;
  assign _01924_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9424" *) mux_265_nl;
  assign _01925_ = or_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9433" *) main_stage_v_4;
  assign _01926_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9433" *) _03900_;
  assign _01927_ = reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9490" *) { lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3] };
  assign _01928_ = _01927_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9490" *) { _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_, _02491_ };
  assign _01929_ = _01928_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9491" *) { _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_, _02591_ };
  assign _01930_ = lut_lookup_if_else_else_else_else_mux_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9494" *) { lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2, lut_lookup_if_else_else_else_asn_mdf_1_sva_2 };
  assign _01931_ = _01930_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9494" *) { _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_, _02592_ };
  assign _01932_ = _01931_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9495" *) { lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8, lut_lookup_1_if_else_slc_32_svs_8 };
  assign _01933_ = lut_lookup_1_else_else_else_else_rshift_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9498" *) { lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4, lut_lookup_else_else_else_asn_mdf_1_sva_4 };
  assign _01934_ = _01933_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9498" *) { lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8, lut_lookup_else_else_slc_32_mdf_1_sva_8 };
  assign _01935_ = lut_lookup_1_else_1_else_else_rshift_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9501" *) { _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_, _02593_ };
  assign _01936_ = _01935_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9501" *) { lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8, lut_lookup_else_1_slc_32_mdf_1_sva_8 };
  assign _01937_ = reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9505" *) { lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3] };
  assign _01938_ = _01937_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9505" *) { _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_, _02493_ };
  assign _01939_ = _01938_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9506" *) { _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_, _02594_ };
  assign _01940_ = lut_lookup_if_else_else_else_else_mux_1_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9509" *) { lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2, lut_lookup_if_else_else_else_asn_mdf_2_sva_2 };
  assign _01941_ = _01940_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9509" *) { _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_, _02595_ };
  assign _01942_ = _01941_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9510" *) { lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8, lut_lookup_2_if_else_slc_32_svs_8 };
  assign _01943_ = lut_lookup_2_else_else_else_else_rshift_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9513" *) { lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4, lut_lookup_else_else_else_asn_mdf_2_sva_4 };
  assign _01944_ = _01943_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9513" *) { lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8, lut_lookup_else_else_slc_32_mdf_2_sva_8 };
  assign _01945_ = lut_lookup_2_else_1_else_else_rshift_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9516" *) { _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_, _02596_ };
  assign _01946_ = _01945_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9516" *) { lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8, lut_lookup_else_1_slc_32_mdf_2_sva_8 };
  assign _01947_ = reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9519" *) { lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3] };
  assign _01948_ = _01947_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9519" *) { _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_, _02495_ };
  assign _01949_ = _01948_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9520" *) { _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_, _02597_ };
  assign _01950_ = lut_lookup_if_else_else_else_else_mux_2_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9523" *) { lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2, lut_lookup_if_else_else_else_asn_mdf_3_sva_2 };
  assign _01951_ = _01950_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9523" *) { _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_, _02598_ };
  assign _01952_ = _01951_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9524" *) { lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8, lut_lookup_3_if_else_slc_32_svs_8 };
  assign _01953_ = lut_lookup_3_else_else_else_else_rshift_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9527" *) { lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4, lut_lookup_else_else_else_asn_mdf_3_sva_4 };
  assign _01954_ = _01953_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9527" *) { lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8, lut_lookup_else_else_slc_32_mdf_3_sva_8 };
  assign _01955_ = lut_lookup_3_else_1_else_else_rshift_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9530" *) { _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_, _02599_ };
  assign _01956_ = _01955_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9530" *) { lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8, lut_lookup_else_1_slc_32_mdf_3_sva_8 };
  assign _01957_ = reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9533" *) { lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3] };
  assign _01958_ = _01957_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9533" *) { _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_, _02497_ };
  assign _01959_ = _01958_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9534" *) { _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_, _02600_ };
  assign _01960_ = lut_lookup_if_else_else_else_else_mux_3_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9537" *) { lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2, lut_lookup_if_else_else_else_asn_mdf_sva_2 };
  assign _01961_ = _01960_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9537" *) { _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_, _02601_ };
  assign _01962_ = _01961_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9538" *) { lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8, lut_lookup_4_if_else_slc_32_svs_8 };
  assign _01963_ = lut_lookup_4_else_else_else_else_rshift_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9541" *) { lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4, lut_lookup_else_else_else_asn_mdf_sva_4 };
  assign _01964_ = _01963_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9541" *) { lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8, lut_lookup_else_else_slc_32_mdf_sva_8 };
  assign _01965_ = lut_lookup_4_else_1_else_else_rshift_itm & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9544" *) { _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_, _02602_ };
  assign _01966_ = _01965_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9544" *) { lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8, lut_lookup_else_1_slc_32_mdf_sva_8 };
  assign _01967_ = lut_lookup_else_mux_180_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9546" *) lut_lookup_lo_uflow_1_lpi_1_dfm_3;
  assign _01968_ = lut_lookup_else_mux_182_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9547" *) lut_lookup_lo_uflow_2_lpi_1_dfm_3;
  assign _01969_ = lut_lookup_else_mux_184_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9548" *) lut_lookup_lo_uflow_3_lpi_1_dfm_3;
  assign _01970_ = lut_lookup_else_mux_186_cse & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9550" *) lut_lookup_lo_uflow_lpi_1_dfm_3;
  assign _01971_ = lut_lookup_if_if_else_else_le_index_s_sva[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9553" *) { lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3], lut_lookup_4_if_if_else_else_if_acc_nl[3] };
  assign _01972_ = _01971_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9553" *) { _02497_, _02497_, _02497_, _02497_, _02497_, _02497_ };
  assign _01973_ = _01972_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9554" *) { _02600_, _02600_, _02600_, _02600_, _02600_, _02600_ };
  assign _01974_ = lut_lookup_if_if_else_else_le_index_s_3_sva[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9562" *) { lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3], lut_lookup_3_if_if_else_else_if_acc_nl[3] };
  assign _01975_ = _01974_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9562" *) { _02495_, _02495_, _02495_, _02495_, _02495_, _02495_ };
  assign _01976_ = _01975_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9563" *) { _02597_, _02597_, _02597_, _02597_, _02597_, _02597_ };
  assign _01977_ = lut_lookup_if_if_else_else_le_index_s_1_sva[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9568" *) { lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3], lut_lookup_1_if_if_else_else_if_acc_nl[3] };
  assign _01978_ = _01977_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9568" *) { _02491_, _02491_, _02491_, _02491_, _02491_, _02491_ };
  assign _01979_ = _01978_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9569" *) { _02591_, _02591_, _02591_, _02591_, _02591_, _02591_ };
  assign _01980_ = lut_lookup_if_if_else_else_le_index_s_2_sva[5:0] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9574" *) { lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3], lut_lookup_2_if_if_else_else_if_acc_nl[3] };
  assign _01981_ = _01980_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9574" *) { _02493_, _02493_, _02493_, _02493_, _02493_, _02493_ };
  assign _01982_ = _01981_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9575" *) { _02594_, _02594_, _02594_, _02594_, _02594_, _02594_ };
  assign _01983_ = mux_1139_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9589" *) or_cse;
  assign _01984_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9590" *) _03901_;
  assign _01985_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9599" *) mux_267_nl;
  assign _01986_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9608" *) mux_268_nl;
  assign _01987_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9617" *) _02603_;
  assign _01988_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9625" *) mux_270_nl;
  assign _01989_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9633" *) _02604_;
  assign _01990_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9653" *) mux_276_nl;
  assign _01991_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9661" *) mux_277_nl;
  assign _01992_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9670" *) mux_278_nl;
  assign _01993_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9679" *) mux_279_nl;
  assign _01994_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9687" *) _02605_;
  assign _01995_ = mux_1152_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9719" *) or_cse;
  assign _01996_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9720" *) _03902_;
  assign _01997_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9729" *) mux_286_nl;
  assign _01998_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9738" *) mux_287_nl;
  assign _01999_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9747" *) mux_289_nl;
  assign _02000_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9755" *) mux_291_nl;
  assign _02001_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9763" *) _02606_;
  assign _02002_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9771" *) _02607_;
  assign _02003_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9779" *) mux_299_nl;
  assign _02004_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9788" *) mux_300_nl;
  assign _02005_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9797" *) _02608_;
  assign _02006_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9805" *) _02609_;
  assign _02007_ = mux_1165_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9813" *) or_cse;
  assign _02008_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9814" *) _03903_;
  assign _02009_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9823" *) mux_308_nl;
  assign _02010_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9832" *) mux_309_nl;
  assign _02011_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9841" *) _02610_;
  assign _02012_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9849" *) mux_311_nl;
  assign _02013_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9867" *) mux_319_nl;
  assign _02014_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9876" *) _02611_;
  assign _02015_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9885" *) _02612_;
  assign _02016_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9893" *) _02613_;
  assign _02017_ = mux_1178_nl & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9911" *) or_cse;
  assign _02018_ = core_wen & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9912" *) _03904_;
  assign _02019_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9921" *) mux_332_nl;
  assign _02020_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9930" *) mux_333_nl;
  assign _02021_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9939" *) _02614_;
  assign _02022_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9947" *) mux_335_nl;
  assign _02023_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9955" *) mux_343_nl;
  assign _02024_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9964" *) _02615_;
  assign _02025_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9973" *) _02616_;
  assign _02026_ = _00924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9981" *) _02617_;
  assign and_dcpl_98 = reg_cfg_precision_1_sva_st_13_cse_1 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12271" *) 2'b10;
  assign _02031_ = chn_lut_in_rsci_d_mxwt[30:23] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13078" *) 8'b11111111;
  assign and_dcpl_309 = cfg_precision_rsci_d == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13115" *) 2'b10;
  assign _02032_ = chn_lut_in_rsci_d_mxwt[126:119] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13120" *) 8'b11111111;
  assign and_956_cse = reg_cfg_precision_1_sva_st_12_cse_1 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5482" *) 2'b10;
  assign and_896_cse = cfg_precision_1_sva_st_70 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5917" *) 2'b10;
  assign _02033_ = FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5962" *) 8'b11111111;
  assign _02034_ = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_2_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6010" *) 8'b11111111;
  assign _02035_ = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_5_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6057" *) 8'b11111111;
  assign _02036_ = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_8_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6097" *) 8'b11111111;
  assign _02037_ = FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_11_tmp == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6138" *) 8'b11111111;
  assign _02038_ = cfg_lut_le_start_rsci_d[30:23] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6153" *) 8'b11111111;
  assign _02039_ = cfg_lut_lo_start_rsci_d[30:23] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6154" *) 8'b11111111;
  assign _02040_ = chn_lut_in_rsci_d_mxwt[62:55] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6155" *) 8'b11111111;
  assign _02041_ = chn_lut_in_rsci_d_mxwt[94:87] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6156" *) 8'b11111111;
  assign lut_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = chn_lut_in_rsci_d_mxwt[30:23] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6176" *) cfg_lut_le_start_rsci_d[30:23];
  assign lut_lookup_1_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp = chn_lut_in_rsci_d_mxwt[30:23] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6178" *) cfg_lut_lo_start_rsci_d[30:23];
  assign lut_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = chn_lut_in_rsci_d_mxwt[62:55] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6180" *) cfg_lut_le_start_rsci_d[30:23];
  assign lut_lookup_2_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp = chn_lut_in_rsci_d_mxwt[62:55] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6182" *) cfg_lut_lo_start_rsci_d[30:23];
  assign lut_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = chn_lut_in_rsci_d_mxwt[94:87] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6184" *) cfg_lut_le_start_rsci_d[30:23];
  assign lut_lookup_3_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp = chn_lut_in_rsci_d_mxwt[94:87] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6186" *) cfg_lut_lo_start_rsci_d[30:23];
  assign lut_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = chn_lut_in_rsci_d_mxwt[126:119] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6188" *) cfg_lut_le_start_rsci_d[30:23];
  assign lut_lookup_4_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp = chn_lut_in_rsci_d_mxwt[126:119] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6190" *) cfg_lut_lo_start_rsci_d[30:23];
  assign _02042_ = FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6216" *) 24'b111111111111111111111111;
  assign _02043_ = FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6232" *) 24'b111111111111111111111111;
  assign _02044_ = FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6256" *) 24'b111111111111111111111111;
  assign _02045_ = FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6272" *) 24'b111111111111111111111111;
  assign _02046_ = FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6296" *) 24'b111111111111111111111111;
  assign _02047_ = FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6312" *) 24'b111111111111111111111111;
  assign _02048_ = FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6336" *) 24'b111111111111111111111111;
  assign _02049_ = FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[48:25] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6352" *) 24'b111111111111111111111111;
  assign _02050_ = cfg_precision_1_sva_8 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6414" *) 2'b10;
  assign _02051_ = FpAdd_8U_23U_o_expo_lpi_1_dfm_7 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6475" *) 8'b11111111;
  assign _02052_ = FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6481" *) 8'b11111111;
  assign _02053_ = FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6662" *) 8'b11111111;
  assign _02054_ = cfg_precision_1_sva_st_71 == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7541" *) 2'b10;
  assign _02055_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10222" *) cfg_lut_lo_start_rsci_d[30:0];
  assign or_1857_cse = cfg_precision_1_sva_st_70 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12053" *) 2'b10;
  assign or_66_cse = reg_cfg_precision_1_sva_st_13_cse_1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12082" *) 2'b10;
  assign or_tmp_314 = cfg_precision_1_sva_st_71 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12377" *) 2'b10;
  assign _02056_ = cfg_precision_1_sva_st_72 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12380" *) 2'b10;
  assign _02057_ = cfg_precision_1_sva_st_107 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12405" *) 2'b10;
  assign or_1202_cse = cfg_precision_1_sva_8 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12962" *) 2'b10;
  assign or_1495_cse = cfg_precision_rsci_d != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13064" *) 2'b10;
  assign or_26_cse = reg_cfg_precision_1_sva_st_12_cse_1 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13067" *) 2'b10;
  assign _02058_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5961" *) FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0;
  assign _02059_ = FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5964" *) 8'b11111111;
  assign _02060_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6009" *) FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_2_mx0;
  assign _02061_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6056" *) FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_2_mx0;
  assign _02062_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6096" *) FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_2_mx0;
  assign _02063_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6137" *) FpAdd_8U_23U_2_o_mant_lpi_1_dfm_2_mx0;
  assign _02064_ = chn_lut_in_rsci_d_mxwt[30:23] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6191" *) 8'b11111111;
  assign _02065_ = chn_lut_in_rsci_d_mxwt[126:119] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6192" *) 8'b11111111;
  assign _02066_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6368" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_2_tmp;
  assign _02067_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6381" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_5_tmp;
  assign _02068_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6396" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_8_tmp;
  assign _02069_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6411" *) FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_11_tmp;
  assign lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6439" *) cfg_lut_le_start_rsci_d[30:0];
  assign lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6440" *) chn_lut_in_rsci_d_mxwt[30:0];
  assign lut_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6445" *) chn_lut_in_rsci_d_mxwt[62:32];
  assign lut_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6450" *) chn_lut_in_rsci_d_mxwt[94:64];
  assign lut_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6455" *) chn_lut_in_rsci_d_mxwt[126:96];
  assign _02070_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6474" *) FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0;
  assign _02071_ = FpAdd_8U_23U_o_expo_lpi_1_dfm_7 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6477" *) 8'b11111111;
  assign _02072_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6480" *) FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0;
  assign _02073_ = FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6483" *) 8'b11111111;
  assign _02074_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6485" *) FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0;
  assign _02075_ = FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7 != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6486" *) 8'b11111111;
  assign _02076_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6550" *) cfg_lut_le_start_rsci_d[22:0];
  assign _02077_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6552" *) cfg_lut_lo_start_rsci_d[22:0];
  assign lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7224" *) lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[286:136];
  assign lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7231" *) lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[286:136];
  assign lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7241" *) lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[286:136];
  assign lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7248" *) lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[286:136];
  assign lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7258" *) lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[286:136];
  assign lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7265" *) lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[286:136];
  assign lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7275" *) lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[286:136];
  assign lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7282" *) lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[286:136];
  assign _02078_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7325" *) chn_lut_in_rsci_d_mxwt[54:32];
  assign _02079_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7326" *) chn_lut_in_rsci_d_mxwt[118:96];
  assign _02080_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7331" *) chn_lut_in_rsci_d_mxwt[22:0];
  assign _02081_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7336" *) chn_lut_in_rsci_d_mxwt[86:64];
  assign _02082_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7379" *) FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:0];
  assign _02083_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7385" *) FpAdd_8U_23U_2_int_mant_p1_1_sva_3[48:0];
  assign _02084_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7391" *) FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:0];
  assign _02085_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7397" *) FpAdd_8U_23U_2_int_mant_p1_2_sva_3[48:0];
  assign _02086_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7403" *) FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:0];
  assign _02087_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7409" *) FpAdd_8U_23U_2_int_mant_p1_3_sva_3[48:0];
  assign _02088_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7415" *) FpAdd_8U_23U_1_int_mant_p1_sva_3[48:0];
  assign _02089_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7421" *) FpAdd_8U_23U_2_int_mant_p1_sva_3[48:0];
  assign _02090_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7456" *) FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp;
  assign _02091_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7458" *) FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7;
  assign _02092_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7460" *) FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7;
  assign _02093_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7462" *) FpAdd_8U_23U_o_expo_lpi_1_dfm_7;
  assign _02094_ = chn_lut_in_rsci_d_mxwt[94:87] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8197" *) 8'b11111111;
  assign _02095_ = chn_lut_in_rsci_d_mxwt[62:55] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8211" *) 8'b11111111;
  assign _02096_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10072" *) lut_lookup_else_1_slc_32_mdf_1_sva_7;
  assign _02097_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10074" *) lut_lookup_else_1_slc_32_mdf_2_sva_7;
  assign _02098_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10076" *) lut_lookup_else_1_slc_32_mdf_3_sva_7;
  assign _02099_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10078" *) lut_lookup_else_1_slc_32_mdf_sva_7;
  assign _02100_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10108" *) mux_tmp_4;
  assign _02101_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10204" *) and_dcpl_54;
  assign _02102_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10204" *) mux_582_itm;
  assign _02103_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10230" *) mux_595_itm;
  assign _02104_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10310" *) cfg_lut_le_start_1_sva_41[31];
  assign _02105_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10319" *) mux_606_nl;
  assign _02106_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10321" *) cfg_lut_lo_start_1_sva_41[31];
  assign _02107_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10330" *) mux_25_itm;
  assign _02108_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10341" *) mux_622_nl;
  assign _02109_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10363" *) mux_634_nl;
  assign _02110_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10385" *) mux_651_nl;
  assign _02111_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10526" *) mux_704_nl;
  assign _02112_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10670" *) cfg_lut_le_function_1_sva_st_41;
  assign _02113_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10671" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
  assign _02114_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10673" *) _02638_;
  assign _02115_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10744" *) lut_lookup_1_if_else_else_else_else_acc_nl[32];
  assign _02116_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10790" *) mux_798_nl;
  assign _02117_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10799" *) mux_799_nl;
  assign _02118_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10808" *) FpAdd_8U_23U_2_mux_13_itm_3;
  assign _02119_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10809" *) FpMantRNE_49U_24U_2_else_carry_1_sva_2;
  assign _02120_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10818" *) mux_1248_nl;
  assign _02121_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10892" *) lut_lookup_2_if_else_else_else_else_acc_nl[32];
  assign _02122_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10922" *) mux_854_nl;
  assign _02123_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10931" *) mux_855_nl;
  assign _02124_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10940" *) FpAdd_8U_23U_2_mux_29_itm_3;
  assign _02125_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10941" *) FpMantRNE_49U_24U_2_else_carry_2_sva_2;
  assign _02126_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10950" *) mux_1250_nl;
  assign _02127_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11012" *) lut_lookup_3_if_else_else_else_else_acc_nl[32];
  assign _02128_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11030" *) mux_910_nl;
  assign _02129_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11039" *) mux_912_nl;
  assign _02130_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11048" *) FpAdd_8U_23U_2_mux_45_itm_3;
  assign _02131_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11049" *) FpMantRNE_49U_24U_2_else_carry_3_sva_2;
  assign _02132_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11138" *) lut_lookup_4_if_else_else_else_else_acc_nl[32];
  assign _02133_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11156" *) mux_969_nl;
  assign _02134_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11165" *) mux_971_nl;
  assign _02135_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11174" *) FpAdd_8U_23U_2_mux_61_itm_3;
  assign _02136_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11175" *) FpMantRNE_49U_24U_2_else_carry_sva_2;
  assign _02137_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11206" *) lut_lookup_else_else_slc_32_mdf_sva_7;
  assign _02138_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11208" *) lut_lookup_else_else_slc_32_mdf_3_sva_7;
  assign _02139_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11210" *) lut_lookup_else_else_slc_32_mdf_2_sva_7;
  assign _02140_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11219" *) lut_lookup_else_else_slc_32_mdf_1_sva_7;
  assign _02141_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11350" *) lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8];
  assign _02142_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11353" *) lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8];
  assign _02143_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11356" *) lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8];
  assign _02144_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11359" *) lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8];
  assign _02145_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11377" *) cfg_lut_le_start_rsci_d[31];
  assign _02146_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11404" *) cfg_lut_lo_start_rsci_d[31];
  assign _02147_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11523" *) mux_1079_nl;
  assign _02148_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11551" *) mux_1086_nl;
  assign _02149_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11579" *) mux_1093_nl;
  assign _02150_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11607" *) mux_1098_nl;
  assign _02151_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11615" *) mux_1101_nl;
  assign _00071_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11747" *) lut_lookup_else_if_lor_5_lpi_1_dfm_6;
  assign _00076_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11750" *) lut_lookup_else_if_lor_6_lpi_1_dfm_6;
  assign _00081_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11753" *) lut_lookup_else_if_lor_7_lpi_1_dfm_6;
  assign _00086_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11756" *) lut_lookup_else_if_lor_1_lpi_1_dfm_6;
  assign _02152_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11759" *) lut_lookup_1_else_2_and_svs;
  assign _02153_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11800" *) lut_lookup_2_else_2_and_svs;
  assign _02154_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11841" *) lut_lookup_3_else_2_and_svs;
  assign _02155_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11882" *) lut_lookup_4_else_2_and_svs;
  assign _00040_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11923" *) chn_lut_in_rsci_d_mxwt[30:23];
  assign _00041_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11924" *) cfg_lut_lo_start_rsci_d[30:23];
  assign _00042_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11930" *) chn_lut_in_rsci_d_mxwt[62:55];
  assign _00043_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11931" *) cfg_lut_le_start_rsci_d[30:23];
  assign _00044_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11937" *) chn_lut_in_rsci_d_mxwt[94:87];
  assign _00045_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11944" *) chn_lut_in_rsci_d_mxwt[126:119];
  assign _02156_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11949" *) FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0;
  assign _02157_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11955" *) FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0;
  assign _02158_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11964" *) FpAdd_8U_23U_2_addend_smaller_qr_1_lpi_1_dfm_mx0;
  assign _02159_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11967" *) FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0;
  assign _02160_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11973" *) FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0;
  assign _02161_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11982" *) FpAdd_8U_23U_2_addend_smaller_qr_2_lpi_1_dfm_mx0;
  assign _02162_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11985" *) FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0;
  assign _02163_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11991" *) FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0;
  assign _02164_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12000" *) FpAdd_8U_23U_2_addend_smaller_qr_3_lpi_1_dfm_mx0;
  assign _02165_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12003" *) FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0;
  assign _02166_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12009" *) FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0;
  assign _02167_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12018" *) FpAdd_8U_23U_2_addend_smaller_qr_lpi_1_dfm_mx0;
  assign _00000_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12021" *) main_stage_v_2;
  assign _00001_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12023" *) main_stage_v_3;
  assign _02168_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12028" *) lut_lookup_1_if_else_slc_32_svs_7;
  assign _02169_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12031" *) FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6;
  assign _02170_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12038" *) mux_1125_nl;
  assign _02171_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12040" *) _01145_;
  assign _00002_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12041" *) or_1936_cse;
  assign _00003_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12045" *) or_1689_cse;
  assign _00004_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12047" *) or_tmp_63;
  assign nor_772_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12050" *) _02654_;
  assign nor_773_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12053" *) _02659_;
  assign nor_769_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12056" *) _02663_;
  assign nor_770_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12060" *) _02666_;
  assign _02172_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12066" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13;
  assign _02173_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12091" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _02174_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12098" *) lut_lookup_2_if_else_slc_32_svs_7;
  assign _02175_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12101" *) FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6;
  assign _02176_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12107" *) mux_1126_cse;
  assign nor_852_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12108" *) _02673_;
  assign nor_760_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12118" *) _02678_;
  assign nor_761_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12121" *) _02682_;
  assign nor_757_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12124" *) _02686_;
  assign nor_758_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12128" *) _02689_;
  assign _02177_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12134" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15;
  assign _02178_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12144" *) _02690_;
  assign _00005_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12148" *) or_tmp_44;
  assign _02179_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12157" *) lut_lookup_3_if_else_slc_32_svs_7;
  assign _02180_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12160" *) FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6;
  assign _02181_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12170" *) _01146_;
  assign _00006_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12171" *) or_tmp_1692;
  assign nor_745_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12180" *) _02698_;
  assign nor_746_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12183" *) _02703_;
  assign nor_742_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12186" *) _02707_;
  assign nor_743_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12190" *) _02710_;
  assign _02182_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12196" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_17;
  assign _02183_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12222" *) lut_lookup_4_if_else_slc_32_svs_7;
  assign _02184_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12225" *) FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6;
  assign _02185_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12235" *) _01147_;
  assign _00007_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12236" *) or_tmp_1705;
  assign nor_732_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12246" *) _02722_;
  assign nor_733_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12249" *) _02726_;
  assign nor_729_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12252" *) _02730_;
  assign nor_730_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12256" *) _02733_;
  assign _02186_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12262" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_19;
  assign nand_76_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12271" *) _01149_;
  assign _02187_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12273" *) or_856_nl;
  assign _02188_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12274" *) _02734_;
  assign _02189_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12280" *) lut_lookup_1_if_else_else_else_if_acc_nl[3];
  assign _02190_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12281" *) and_tmp_5;
  assign _02191_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12283" *) lut_lookup_else_else_else_asn_mdf_1_sva_st_3;
  assign nor_726_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12287" *) _02738_;
  assign nor_727_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12288" *) _02739_;
  assign nor_881_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12290" *) _02740_;
  assign nor_721_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12293" *) _02741_;
  assign _02192_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12301" *) lut_lookup_2_if_else_else_else_if_acc_nl[3];
  assign _02193_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12302" *) and_tmp_27;
  assign _02194_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12304" *) lut_lookup_else_else_else_asn_mdf_2_sva_st_3;
  assign nor_719_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12308" *) _02744_;
  assign nor_720_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12309" *) _02745_;
  assign nor_713_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12311" *) _02746_;
  assign nor_714_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12314" *) _02747_;
  assign _02195_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12322" *) lut_lookup_3_if_else_else_else_if_acc_nl[3];
  assign _02196_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12323" *) and_tmp_14;
  assign nor_711_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12328" *) _02749_;
  assign nor_712_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12329" *) _02750_;
  assign nor_880_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12331" *) _02751_;
  assign _00008_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12334" *) or_tmp_378;
  assign _02197_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12341" *) lut_lookup_4_if_else_else_else_if_acc_nl[3];
  assign _02198_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12342" *) and_tmp_19;
  assign _02199_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12344" *) lut_lookup_else_else_else_asn_mdf_sva_st_3;
  assign nor_705_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12348" *) _02754_;
  assign nor_706_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12349" *) _02755_;
  assign nor_879_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12351" *) _02756_;
  assign nor_700_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12354" *) _02757_;
  assign _00009_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12370" *) mux_tmp_1136;
  assign _02200_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12374" *) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9];
  assign _02201_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12375" *) cfg_lut_le_function_1_sva_st_42;
  assign _00032_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12377" *) main_stage_v_4;
  assign nor_698_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12377" *) _02763_;
  assign _02202_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12378" *) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  assign _02203_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12380" *) and_843_cse;
  assign nor_699_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12380" *) _02768_;
  assign nor_696_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12384" *) _02772_;
  assign nor_697_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12386" *) _02775_;
  assign nor_694_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12393" *) _02782_;
  assign nor_695_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12394" *) _02783_;
  assign _00010_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12396" *) main_stage_v_5;
  assign _02204_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12400" *) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9];
  assign nor_692_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12402" *) _02787_;
  assign _02205_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12403" *) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  assign nor_693_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12406" *) _02792_;
  assign nor_691_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12409" *) _02795_;
  assign nor_689_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12412" *) _02798_;
  assign _00011_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12417" *) mux_tmp_1149;
  assign _02206_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12421" *) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9];
  assign nor_686_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12424" *) _02807_;
  assign _02207_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12425" *) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  assign nor_687_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12427" *) _02812_;
  assign nor_684_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12430" *) _02816_;
  assign nor_685_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12432" *) _02819_;
  assign nor_681_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12436" *) _02823_;
  assign _02208_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12437" *) cfg_lut_le_function_1_sva_10;
  assign nor_682_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12438" *) _02826_;
  assign nor_683_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12440" *) _02829_;
  assign nor_678_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12445" *) _02831_;
  assign nor_679_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12448" *) _02832_;
  assign nor_680_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12450" *) _02833_;
  assign _02209_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12457" *) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9];
  assign nor_676_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12459" *) _02837_;
  assign _02210_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12460" *) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  assign nor_677_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12462" *) _02842_;
  assign nor_674_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12465" *) or_365_cse;
  assign nor_675_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12467" *) _02846_;
  assign _00012_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12472" *) mux_tmp_1162;
  assign _02211_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12476" *) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9];
  assign nor_672_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12479" *) _02852_;
  assign _02212_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12480" *) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  assign nor_673_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12482" *) _02857_;
  assign nor_670_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12486" *) _02861_;
  assign nor_671_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12488" *) _02864_;
  assign nor_668_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12495" *) _02871_;
  assign nor_669_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12496" *) _02872_;
  assign _02213_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12498" *) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9];
  assign nor_666_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12500" *) _02876_;
  assign _02214_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12501" *) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  assign nor_667_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12504" *) _02881_;
  assign _00013_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12515" *) mux_tmp_1175;
  assign _02215_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12519" *) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9];
  assign nor_664_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12522" *) _02894_;
  assign _02216_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12523" *) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  assign nor_665_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12525" *) _02899_;
  assign nor_662_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12529" *) _02903_;
  assign nor_663_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12531" *) _02906_;
  assign nor_660_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12538" *) _02913_;
  assign nor_661_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12539" *) _02914_;
  assign _02217_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12541" *) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9];
  assign nor_658_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12543" *) _02918_;
  assign _02218_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12544" *) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  assign nor_659_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12546" *) _02923_;
  assign _02219_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12557" *) lut_lookup_else_else_else_asn_mdf_sva_4;
  assign _02220_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12560" *) _02931_;
  assign lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_4_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12562" *) _02933_;
  assign _02221_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12563" *) lut_lookup_else_else_else_asn_mdf_3_sva_4;
  assign _02222_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12566" *) _02934_;
  assign lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_5_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12568" *) _02936_;
  assign _02223_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12569" *) lut_lookup_else_else_else_asn_mdf_2_sva_4;
  assign _02224_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12572" *) _02937_;
  assign lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_6_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12574" *) _02939_;
  assign _02225_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12575" *) lut_lookup_else_else_else_asn_mdf_1_sva_4;
  assign _02226_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12578" *) _02940_;
  assign lut_lookup_if_if_lut_lookup_if_if_lut_lookup_if_if_nor_7_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12580" *) _02942_;
  assign _02227_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12612" *) mux_tmp_595;
  assign _00014_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12614" *) mux_598_nl;
  assign _02228_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12621" *) or_186_nl;
  assign _02229_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12622" *) reg_chn_lut_out_rsci_ld_core_psct_cse;
  assign _00015_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12624" *) mux_611_nl;
  assign _02230_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12628" *) mux_477_nl;
  assign nand_15_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12628" *) _01164_;
  assign nand_16_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12637" *) _01165_;
  assign _02231_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12643" *) mux_534_nl;
  assign nand_17_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12643" *) _01166_;
  assign _02232_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12651" *) and_tmp_59;
  assign nor_642_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12651" *) _02945_;
  assign _02233_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12692" *) _02947_;
  assign nor_792_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12693" *) or_1857_cse;
  assign nor_638_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12693" *) _02948_;
  assign _00017_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12697" *) mux_662_nl;
  assign _02234_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12699" *) _02950_;
  assign _02235_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12701" *) lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02236_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12704" *) or_tmp_314;
  assign nor_640_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12704" *) _02951_;
  assign _02237_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12705" *) lut_lookup_4_if_else_slc_32_svs_st_5;
  assign _02238_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12706" *) lut_lookup_if_else_else_else_asn_mdf_sva_2;
  assign _00018_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12708" *) mux_665_nl;
  assign _02239_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12713" *) _02955_;
  assign nor_633_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12714" *) _02956_;
  assign _00019_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12718" *) mux_673_nl;
  assign nand_18_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12720" *) _01181_;
  assign nor_636_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12722" *) _02958_;
  assign _02240_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12723" *) lut_lookup_3_if_else_slc_32_svs_st_5;
  assign _02241_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12724" *) lut_lookup_if_else_else_else_asn_mdf_3_sva_2;
  assign _00020_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12726" *) mux_676_nl;
  assign _02242_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12730" *) _02962_;
  assign nor_628_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12731" *) _02963_;
  assign _00021_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12735" *) mux_684_nl;
  assign nand_19_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12737" *) _01182_;
  assign nor_631_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12739" *) _02965_;
  assign _02243_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12740" *) lut_lookup_2_if_else_slc_32_svs_st_5;
  assign _02244_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12741" *) lut_lookup_if_else_else_else_asn_mdf_2_sva_2;
  assign _00022_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12743" *) mux_687_nl;
  assign _02245_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12746" *) lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1;
  assign nor_623_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12747" *) _02968_;
  assign _00023_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12751" *) mux_695_nl;
  assign _02246_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12753" *) lut_lookup_else_unequal_tmp_18;
  assign _02247_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12754" *) _02970_;
  assign nand_20_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12754" *) _01183_;
  assign nor_626_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12756" *) _02971_;
  assign _02248_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12757" *) lut_lookup_1_if_else_slc_32_svs_st_5;
  assign _02249_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12758" *) lut_lookup_if_else_else_else_asn_mdf_1_sva_2;
  assign _00024_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12760" *) mux_698_nl;
  assign _02250_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12764" *) _02975_;
  assign _02251_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12768" *) _02978_;
  assign nor_619_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12773" *) _02981_;
  assign _02252_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12782" *) _01184_;
  assign nor_616_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12782" *) _02984_;
  assign _00025_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12785" *) mux_755_cse;
  assign _00026_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12790" *) mux_758_nl;
  assign _00027_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12796" *) or_tmp_993;
  assign nor_831_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12801" *) _02986_;
  assign nor_833_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12804" *) _02988_;
  assign nor_597_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12809" *) _02994_;
  assign _02253_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12810" *) IsNaN_8U_23U_6_land_1_lpi_1_dfm_6;
  assign _02254_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12811" *) lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02255_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12815" *) _01187_;
  assign nor_598_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12815" *) _03001_;
  assign _02256_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12824" *) nor_tmp_238;
  assign nor_595_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12824" *) _03002_;
  assign _02257_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12833" *) and_tmp_98;
  assign _02258_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12835" *) FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5;
  assign _02259_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12837" *) or_tmp_1716;
  assign nor_830_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12837" *) _03006_;
  assign _00028_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12850" *) mux_822_nl;
  assign _02260_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12862" *) _01195_;
  assign nor_575_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12862" *) _03011_;
  assign _02261_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *) _01200_;
  assign nor_576_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *) _03016_;
  assign _02262_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12873" *) nor_tmp_260;
  assign nor_573_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12873" *) _03017_;
  assign _02263_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12880" *) and_tmp_108;
  assign _02264_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12882" *) FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5;
  assign _00029_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12897" *) mux_877_nl;
  assign nor_551_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12909" *) _03026_;
  assign _02265_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12910" *) lut_lookup_else_else_else_asn_mdf_3_sva_st_3;
  assign _02266_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *) _01212_;
  assign nor_552_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *) _03031_;
  assign _02267_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12920" *) nor_tmp_281;
  assign nor_549_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12920" *) _03032_;
  assign _02268_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12927" *) and_tmp_119;
  assign _02269_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12929" *) FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5;
  assign nor_827_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12930" *) _03036_;
  assign nand_102_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12932" *) _01218_;
  assign _02270_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12939" *) _01219_;
  assign nor_544_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12939" *) _03039_;
  assign _00030_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12942" *) mux_745_cse;
  assign _02271_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12945" *) _01220_;
  assign nor_540_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12945" *) _03042_;
  assign _00031_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12953" *) mux_935_nl;
  assign nor_528_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12969" *) _03048_;
  assign _02272_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12971" *) IsNaN_8U_23U_6_land_lpi_1_dfm_6;
  assign _02273_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12974" *) _01223_;
  assign nor_529_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12974" *) _03055_;
  assign _02274_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12988" *) and_tmp_131;
  assign _02275_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12990" *) FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5;
  assign nor_825_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12991" *) _03059_;
  assign nand_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12993" *) _01231_;
  assign _02276_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12999" *) _01233_;
  assign nor_518_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12999" *) _03064_;
  assign nor_519_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13001" *) _03067_;
  assign nor_521_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13003" *) or_1931_nl;
  assign _02277_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13016" *) _01235_;
  assign nor_512_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13016" *) _03071_;
  assign nor_513_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13018" *) _03073_;
  assign nor_515_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13020" *) or_1948_nl;
  assign _02278_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13032" *) _01237_;
  assign nor_506_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13032" *) _03077_;
  assign nor_507_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13034" *) _03079_;
  assign nor_509_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13036" *) or_1964_nl;
  assign _02279_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13048" *) _01239_;
  assign nor_500_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13048" *) _03083_;
  assign nor_501_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13050" *) _03085_;
  assign nor_503_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13052" *) or_1983_nl;
  assign _02280_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13065" *) chn_lut_in_rsci_bawt;
  assign nor_495_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13065" *) _03090_;
  assign _02281_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13066" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign _00033_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13066" *) main_stage_v_1;
  assign nor_496_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13067" *) _03093_;
  assign _02282_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13069" *) _03094_;
  assign nor_497_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13070" *) _03097_;
  assign _02283_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13074" *) _01240_;
  assign nor_493_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13074" *) _03099_;
  assign nor_494_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13076" *) _03100_;
  assign nor_491_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13079" *) _03102_;
  assign nor_492_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13081" *) _03104_;
  assign nor_489_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13084" *) _03107_;
  assign nor_490_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13086" *) _03109_;
  assign nor_487_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13088" *) _03110_;
  assign nor_488_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13090" *) _03113_;
  assign nor_485_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13093" *) _03116_;
  assign nor_486_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13095" *) _03118_;
  assign nor_483_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13097" *) _03119_;
  assign nor_484_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13099" *) _03121_;
  assign nor_480_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13102" *) _03124_;
  assign nor_481_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13104" *) _03126_;
  assign nor_475_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13107" *) _03129_;
  assign nor_476_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13109" *) _03130_;
  assign _02284_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13111" *) _03131_;
  assign nor_477_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13112" *) _03134_;
  assign _02285_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13115" *) _01243_;
  assign nor_472_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13116" *) _03135_;
  assign nor_473_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13118" *) _03138_;
  assign nor_470_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13121" *) _03140_;
  assign nor_471_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13123" *) _03142_;
  assign nor_467_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13126" *) _03145_;
  assign nor_468_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13128" *) _03147_;
  assign _02286_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13133" *) lut_lookup_1_if_else_slc_32_svs_6;
  assign _02287_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13134" *) _01248_;
  assign nor_463_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13134" *) _03149_;
  assign nor_464_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13139" *) _03152_;
  assign _02288_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13146" *) lut_lookup_else_1_slc_32_mdf_1_sva_6;
  assign _02289_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13147" *) and_tmp_61;
  assign _02290_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13153" *) and_193_nl;
  assign nor_459_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13153" *) _03154_;
  assign _02291_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13164" *) _01258_;
  assign _02292_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13170" *) and_204_nl;
  assign nor_455_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13170" *) _03155_;
  assign _02293_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13179" *) lut_lookup_else_1_slc_32_mdf_3_sva_6;
  assign _02294_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13180" *) and_tmp_69;
  assign _02295_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13185" *) lut_lookup_4_if_else_slc_32_svs_6;
  assign _02296_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13186" *) _01264_;
  assign nor_453_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13186" *) _03158_;
  assign nor_454_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13190" *) _03161_;
  assign _02297_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13199" *) _01270_;
  assign nand_33_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13201" *) _01271_;
  assign _02298_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13209" *) _01274_;
  assign nor_451_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13209" *) _03162_;
  assign _02299_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13211" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _02300_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13213" *) FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5;
  assign _02301_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13214" *) _01276_;
  assign nor_450_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13214" *) _03165_;
  assign _02302_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13218" *) FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5;
  assign _02303_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13219" *) _01278_;
  assign nor_448_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13219" *) _03168_;
  assign _02304_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13221" *) _01280_;
  assign nor_449_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13221" *) _03169_;
  assign nand_113_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13234" *) _01281_;
  assign _02305_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13236" *) mux_tmp_1247;
  assign nand_114_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13239" *) _01282_;
  assign nand_115_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13247" *) _01283_;
  assign _02306_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13249" *) mux_tmp_1250;
  assign nand_116_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13252" *) _01284_;
  assign nand_117_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13260" *) _01285_;
  assign _02307_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13262" *) mux_tmp_1253;
  assign nand_118_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13265" *) _01286_;
  assign _02308_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13273" *) mux_tmp_1257;
  assign nor_882_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13273" *) _03174_;
  assign _02309_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13276" *) mux_1297_nl;
  assign nl_lut_lookup_1_IntLog2_32U_lshift_rg_s[4:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4391" *) reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[4:0];
  assign nl_lut_lookup_2_IntLog2_32U_lshift_rg_s[4:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4394" *) reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[4:0];
  assign nl_lut_lookup_3_IntLog2_32U_lshift_rg_s[4:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4397" *) reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[4:0];
  assign nl_lut_lookup_4_IntLog2_32U_lshift_rg_s[4:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4400" *) reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[4:0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4422" *) FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm[0];
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4428" *) FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm[0];
  assign _02310_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4447" *) FpAdd_8U_23U_2_b_right_shift_qr_1_lpi_1_dfm[7:1];
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4451" *) FpAdd_8U_23U_2_b_right_shift_qr_1_lpi_1_dfm[0];
  assign _02311_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4458" *) FpAdd_8U_23U_2_a_right_shift_qr_1_lpi_1_dfm[7:1];
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4462" *) FpAdd_8U_23U_2_a_right_shift_qr_1_lpi_1_dfm[0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4468" *) FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm[0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4474" *) FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm[0];
  assign _02312_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4493" *) FpAdd_8U_23U_2_b_right_shift_qr_2_lpi_1_dfm[7:1];
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4497" *) FpAdd_8U_23U_2_b_right_shift_qr_2_lpi_1_dfm[0];
  assign _02313_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4504" *) FpAdd_8U_23U_2_a_right_shift_qr_2_lpi_1_dfm[7:1];
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4508" *) FpAdd_8U_23U_2_a_right_shift_qr_2_lpi_1_dfm[0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4514" *) FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm[0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4520" *) FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm[0];
  assign _02314_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4539" *) FpAdd_8U_23U_2_b_right_shift_qr_3_lpi_1_dfm[7:1];
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4543" *) FpAdd_8U_23U_2_b_right_shift_qr_3_lpi_1_dfm[0];
  assign _02315_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4550" *) FpAdd_8U_23U_2_a_right_shift_qr_3_lpi_1_dfm[7:1];
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4554" *) FpAdd_8U_23U_2_a_right_shift_qr_3_lpi_1_dfm[0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4560" *) FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm[0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4566" *) FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm[0];
  assign _02316_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4585" *) FpAdd_8U_23U_2_b_right_shift_qr_lpi_1_dfm[7:1];
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4589" *) FpAdd_8U_23U_2_b_right_shift_qr_lpi_1_dfm[0];
  assign _02317_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4596" *) FpAdd_8U_23U_2_a_right_shift_qr_lpi_1_dfm[7:1];
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4600" *) FpAdd_8U_23U_2_a_right_shift_qr_lpi_1_dfm[0];
  assign _02318_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5452" *) _03351_;
  assign _02319_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5461" *) lut_lookup_unequal_tmp_13;
  assign _02320_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5471" *) mux_4_nl;
  assign nor_193_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5475" *) or_66_cse;
  assign nor_783_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5475" *) _03356_;
  assign _02321_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5483" *) reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign _02322_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5488" *) mux_20_itm;
  assign nor_874_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5494" *) or_cse;
  assign _02323_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5496" *) _03357_;
  assign _02324_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5501" *) reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign _02325_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5503" *) _03358_;
  assign _02326_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5505" *) mux_26_itm;
  assign _02327_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5510" *) reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign _02328_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5512" *) _03359_;
  assign _02329_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5519" *) reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign nor_775_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5533" *) _03364_;
  assign nor_776_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5536" *) _03369_;
  assign _02330_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5540" *) FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49];
  assign nor_5_cse_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5540" *) _03370_;
  assign _02331_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5542" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12;
  assign _02332_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5550" *) lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7];
  assign _02333_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5556" *) _03372_;
  assign nor_865_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5558" *) _03373_;
  assign _02334_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5562" *) mux_83_cse;
  assign _02335_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5564" *) FpAdd_8U_23U_2_int_mant_p1_1_sva_3[49];
  assign nor_13_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5564" *) _03374_;
  assign FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5568" *) _03375_;
  assign _02336_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5569" *) lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7];
  assign nor_764_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5582" *) _03381_;
  assign nor_765_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5585" *) _03385_;
  assign _02337_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5590" *) FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49];
  assign nor_27_cse_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5590" *) _03386_;
  assign _02338_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5592" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14;
  assign _02339_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5600" *) lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7];
  assign nor_855_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5606" *) _03388_;
  assign _02340_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5611" *) FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49];
  assign nor_31_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5611" *) _03389_;
  assign FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5613" *) _03390_;
  assign _02341_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5614" *) lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7];
  assign _02342_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5619" *) mux_132_nl;
  assign _02343_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5620" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign nor_749_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5623" *) _03395_;
  assign nor_750_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5626" *) _03399_;
  assign _02344_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5630" *) FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49];
  assign nor_38_cse_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5630" *) _03400_;
  assign _02345_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5632" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_16;
  assign _02346_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5640" *) lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7];
  assign _02347_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5644" *) FpAdd_8U_23U_2_int_mant_p1_3_sva_3[49];
  assign nor_42_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5644" *) _03401_;
  assign FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5647" *) _03402_;
  assign _02348_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5648" *) lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7];
  assign nor_737_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5654" *) _03407_;
  assign nor_738_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5657" *) _03411_;
  assign _02349_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5661" *) FpAdd_8U_23U_1_int_mant_p1_sva_3[49];
  assign nor_50_cse_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5661" *) _03412_;
  assign _02350_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5663" *) libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_18;
  assign _02351_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5671" *) lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7];
  assign _02352_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5675" *) FpAdd_8U_23U_2_int_mant_p1_sva_3[49];
  assign nor_54_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5675" *) _03413_;
  assign FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5677" *) _03414_;
  assign _02353_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5678" *) lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7];
  assign _02354_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5687" *) and_tmp_6;
  assign nor_724_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5687" *) _03415_;
  assign _02355_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5688" *) and_tmp_83;
  assign nor_725_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5688" *) _03416_;
  assign nor_722_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5693" *) _03421_;
  assign nor_723_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5695" *) _03424_;
  assign _02356_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5705" *) mux_226_nl;
  assign nor_715_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5708" *) _03430_;
  assign nor_716_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5710" *) _03432_;
  assign _02357_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5717" *) mux_238_nl;
  assign nor_707_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5721" *) _03437_;
  assign nor_708_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5723" *) _03440_;
  assign _02358_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5729" *) mux_251_nl;
  assign nor_701_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5732" *) _03445_;
  assign nor_702_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5734" *) _03448_;
  assign _02359_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5740" *) mux_263_nl;
  assign _02360_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5747" *) mux_275_nl;
  assign nor_690_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5750" *) or_332_nl;
  assign _02361_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5754" *) mux_284_nl;
  assign _02362_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5756" *) mux_285_nl;
  assign _02363_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5768" *) mux_316_nl;
  assign _02364_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5772" *) mux_330_nl;
  assign _02365_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5780" *) and_832_cse;
  assign nor_657_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5780" *) _03450_;
  assign nor_610_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5784" *) or_1202_cse;
  assign _02366_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5801" *) mux_3_itm;
  assign _02367_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5810" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl[23];
  assign _02368_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5813" *) cfg_lut_le_function_rsci_d;
  assign _02369_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5818" *) FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl[23];
  assign _02370_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5822" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl[23];
  assign _02371_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5826" *) FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl[23];
  assign _02372_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5828" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl[23];
  assign _02373_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5830" *) FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl[23];
  assign _02374_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5833" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl[23];
  assign _02375_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5835" *) FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl[23];
  assign _02377_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5853" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _02378_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5856" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
  assign _02379_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5862" *) IsNaN_8U_23U_8_land_2_lpi_1_dfm_5;
  assign nor_190_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5866" *) or_26_cse;
  assign _02380_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5867" *) IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
  assign _02381_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5869" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _02382_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5878" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  assign _02385_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5895" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _02386_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5898" *) reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse;
  assign _02388_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5910" *) mux_671_nl;
  assign _02389_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5912" *) lut_lookup_else_unequal_tmp_12;
  assign nor_634_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5912" *) _03460_;
  assign _02390_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5921" *) mux_717_nl;
  assign _02391_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5925" *) mux_735_nl;
  assign _02392_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5935" *) mux_749_nl;
  assign nor_612_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5938" *) or_978_cse;
  assign nor_606_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5940" *) _03065_;
  assign nor_609_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5944" *) _03462_;
  assign _02393_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5956" *) IsNaN_8U_23U_3_land_1_lpi_1_dfm_6;
  assign _02394_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5963" *) _02058_;
  assign nor_832_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5964" *) _03463_;
  assign nor_434_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5965" *) _03464_;
  assign nor_435_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5966" *) _03465_;
  assign nor_432_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5975" *) _03467_;
  assign nor_433_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5977" *) _03469_;
  assign nor_430_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5980" *) _03470_;
  assign _02395_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5982" *) _01605_;
  assign nor_431_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5982" *) _03471_;
  assign _02396_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6000" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_7;
  assign { _00066_[7], _00066_[5:0] } = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6004" *) cfg_lut_lo_index_select_1_sva_6[7:1];
  assign _02397_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6014" *) _01609_;
  assign nor_588_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6014" *) _03474_;
  assign _02398_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6020" *) IsNaN_8U_23U_3_land_2_lpi_1_dfm_7;
  assign nor_426_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6033" *) _03476_;
  assign nor_427_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6035" *) _03478_;
  assign nor_424_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6038" *) _03479_;
  assign _02399_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6040" *) _01610_;
  assign nor_425_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6040" *) _03480_;
  assign _02400_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6055" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_7;
  assign _02401_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6060" *) _01612_;
  assign nor_564_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6060" *) _03483_;
  assign _02402_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6066" *) IsNaN_8U_23U_3_land_3_lpi_1_dfm_7;
  assign nor_420_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6078" *) _03485_;
  assign nor_421_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6080" *) _03487_;
  assign nor_418_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6083" *) _03488_;
  assign _02403_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6084" *) lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign nor_419_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6085" *) _03490_;
  assign _02404_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6095" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_7;
  assign _02405_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6108" *) IsNaN_8U_23U_3_land_lpi_1_dfm_6;
  assign nor_414_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6120" *) _03492_;
  assign nor_415_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6121" *) _03493_;
  assign nor_412_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6124" *) _03494_;
  assign nor_413_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6125" *) _03495_;
  assign nor_526_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6131" *) _03496_;
  assign _02406_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6136" *) IsNaN_8U_23U_7_land_lpi_1_dfm_7;
  assign nor_482_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6157" *) _02383_;
  assign nor_478_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6158" *) _03498_;
  assign nor_479_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6160" *) _03500_;
  assign nor_469_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6164" *) _02387_;
  assign nor_465_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6166" *) _03501_;
  assign nor_466_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6168" *) _03502_;
  assign IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6191" *) _03503_;
  assign IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6192" *) _03504_;
  assign _00062_[4:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6194" *) reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[4:0];
  assign _00063_[4:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6234" *) reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[4:0];
  assign _00064_[4:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6274" *) reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[4:0];
  assign _00065_[4:0] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6314" *) reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[4:0];
  assign { _00067_[7], _00067_[5:0] } = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6360" *) cfg_lut_le_index_select_1_sva_6[7:1];
  assign IsZero_8U_23U_8_IsZero_8U_23U_8_nor_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6368" *) _03698_;
  assign IsZero_8U_23U_8_IsZero_8U_23U_8_nor_1_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6381" *) _03700_;
  assign IsZero_8U_23U_8_IsZero_8U_23U_8_nor_2_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6396" *) _03702_;
  assign IsZero_8U_23U_8_IsZero_8U_23U_8_nor_3_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6411" *) _03704_;
  assign lut_lookup_if_unequal_tmp_1_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6414" *) _02050_;
  assign _02407_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6416" *) lut_lookup_4_if_else_slc_32_svs_8;
  assign _02408_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6422" *) lut_lookup_3_if_else_slc_32_svs_8;
  assign _02409_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6428" *) lut_lookup_2_if_else_slc_32_svs_8;
  assign _02410_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6434" *) lut_lookup_1_if_else_slc_32_svs_8;
  assign IsNaN_8U_23U_4_land_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6460" *) _02384_;
  assign IsNaN_8U_23U_4_land_1_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6461" *) _02376_;
  assign _02411_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6476" *) _02070_;
  assign _02412_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6477" *) _03705_;
  assign lut_lookup_unequal_tmp_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6479" *) and_896_cse;
  assign _02413_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6482" *) _02072_;
  assign _02414_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6483" *) _03707_;
  assign _02415_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6485" *) _02074_;
  assign _02416_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6486" *) _03709_;
  assign IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6549" *) _03712_;
  assign IsNaN_8U_23U_4_nor_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6550" *) _02076_;
  assign IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6551" *) _02038_;
  assign IsNaN_8U_23U_8_nor_2_tmp_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6552" *) _02077_;
  assign IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_mx0w0 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6553" *) _02039_;
  assign _02417_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6587" *) lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7];
  assign _02418_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6595" *) _03713_;
  assign _02419_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6597" *) FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0;
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6609" *) _03714_;
  assign _02420_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6615" *) lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7];
  assign _02421_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6623" *) _03715_;
  assign _02422_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6625" *) FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_5_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6636" *) _02664_;
  assign _02423_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6638" *) lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7];
  assign _02424_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6646" *) _03716_;
  assign _02425_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6648" *) FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0;
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6660" *) _03717_;
  assign _02426_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6668" *) lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7];
  assign _02427_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6676" *) _03718_;
  assign _02428_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6678" *) FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_7_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6689" *) _02687_;
  assign _02429_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6691" *) lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7];
  assign _02430_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6699" *) _03719_;
  assign _02431_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6701" *) FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0;
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6713" *) _03720_;
  assign _02432_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6719" *) lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7];
  assign _02433_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6727" *) _03721_;
  assign _02434_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6729" *) FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_9_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6740" *) _02708_;
  assign _02435_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6742" *) lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7];
  assign _02436_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6750" *) _03722_;
  assign _02437_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6752" *) FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0;
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6764" *) _03723_;
  assign _02438_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6770" *) lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7];
  assign _02439_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6778" *) _03724_;
  assign _02440_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6780" *) FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_nor_11_m1c = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6791" *) _02731_;
  assign lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6848" *) _03170_;
  assign _00074_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6854" *) lut_lookup_if_1_lor_5_lpi_1_dfm_5;
  assign lut_lookup_1_else_2_else_lut_lookup_else_2_else_if_nor_svs = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6867" *) _03725_;
  assign _00070_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6871" *) IsNaN_8U_23U_6_land_1_lpi_1_dfm_7;
  assign _02441_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6874" *) FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_1_sva_2[255:9];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6877" *) _00046_;
  assign lut_lookup_else_if_else_le_int_1_lpi_1_dfm_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6879" *) _00047_;
  assign _02442_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6881" *) FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2[255:9];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6885" *) _00048_;
  assign lut_lookup_if_1_else_lo_int_1_lpi_1_dfm_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6887" *) _00049_;
  assign _00073_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6889" *) lut_lookup_if_1_else_lo_int_1_lpi_1_dfm_1[8];
  assign _00072_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6894" *) IsNaN_8U_23U_10_land_1_lpi_1_dfm_6;
  assign lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6907" *) _03171_;
  assign _00079_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6913" *) lut_lookup_if_1_lor_6_lpi_1_dfm_5;
  assign lut_lookup_2_else_2_else_lut_lookup_else_2_else_if_nor_svs = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6925" *) _03726_;
  assign _00075_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6929" *) IsNaN_8U_23U_6_land_2_lpi_1_dfm_7;
  assign _02443_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6932" *) FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_2_sva_2[255:9];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6935" *) _00050_;
  assign lut_lookup_else_if_else_le_int_2_lpi_1_dfm_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6937" *) _00051_;
  assign _02444_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6939" *) FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2[255:9];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_1_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6943" *) _00052_;
  assign lut_lookup_if_1_else_lo_int_2_lpi_1_dfm_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6945" *) _00053_;
  assign _00078_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6947" *) lut_lookup_if_1_else_lo_int_2_lpi_1_dfm_1[8];
  assign _00077_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6952" *) IsNaN_8U_23U_10_land_2_lpi_1_dfm_6;
  assign lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6965" *) _03172_;
  assign _00084_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6971" *) lut_lookup_if_1_lor_7_lpi_1_dfm_5;
  assign lut_lookup_3_else_2_else_lut_lookup_else_2_else_if_nor_svs = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6983" *) _03727_;
  assign _00080_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6987" *) IsNaN_8U_23U_6_land_3_lpi_1_dfm_7;
  assign _02445_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6990" *) FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_3_sva_2[255:9];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6993" *) _00054_;
  assign lut_lookup_else_if_else_le_int_3_lpi_1_dfm_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6995" *) _00055_;
  assign _02446_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6997" *) FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2[255:9];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_2_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7001" *) _00056_;
  assign lut_lookup_if_1_else_lo_int_3_lpi_1_dfm_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7003" *) _00057_;
  assign _00083_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7005" *) lut_lookup_if_1_else_lo_int_3_lpi_1_dfm_1[8];
  assign _00082_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7010" *) IsNaN_8U_23U_10_land_3_lpi_1_dfm_6;
  assign _00089_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7021" *) lut_lookup_if_1_lor_1_lpi_1_dfm_5;
  assign lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7029" *) _03173_;
  assign lut_lookup_4_else_2_else_lut_lookup_else_2_else_if_nor_svs = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7041" *) _03728_;
  assign _00085_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7045" *) IsNaN_8U_23U_6_land_lpi_1_dfm_7;
  assign _02447_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7048" *) FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_sva_2[255:9];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7051" *) _00058_;
  assign lut_lookup_else_if_else_le_int_lpi_1_dfm_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7053" *) _00059_;
  assign _02028_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7055" *) FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2[255:9];
  assign FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_3_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7059" *) _00060_;
  assign lut_lookup_if_1_else_lo_int_lpi_1_dfm_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7061" *) _00061_;
  assign _00088_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7063" *) lut_lookup_if_1_else_lo_int_lpi_1_dfm_1[8];
  assign _00087_[34] = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7068" *) IsNaN_8U_23U_10_land_lpi_1_dfm_6;
  assign lut_lookup_lut_lookup_nor_19_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7073" *) lut_lookup_not_39_nl;
  assign _02448_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7075" *) lut_lookup_or_3_tmp;
  assign _02449_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7081" *) _03730_;
  assign _02450_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7084" *) _03732_;
  assign _02451_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7085" *) lut_lookup_1_and_svs_2;
  assign lut_lookup_lut_lookup_nor_18_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7087" *) lut_lookup_not_38_nl;
  assign _02452_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7089" *) lut_lookup_or_7_tmp;
  assign _02453_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7090" *) lut_lookup_else_unequal_tmp_13;
  assign _02454_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7095" *) _03734_;
  assign _02455_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7098" *) _03736_;
  assign _02456_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7099" *) lut_lookup_2_and_svs_2;
  assign lut_lookup_lut_lookup_nor_17_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7101" *) lut_lookup_not_37_nl;
  assign _02457_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7103" *) lut_lookup_or_11_tmp;
  assign _02458_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7109" *) _03738_;
  assign _02459_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7112" *) _03740_;
  assign _02460_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7113" *) lut_lookup_3_and_svs_2;
  assign lut_lookup_lut_lookup_nor_16_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7115" *) lut_lookup_not_36_nl;
  assign _02461_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7117" *) lut_lookup_or_15_tmp;
  assign _02462_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7123" *) _03742_;
  assign _02463_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7126" *) _03744_;
  assign _02464_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7127" *) lut_lookup_4_and_svs_2;
  assign IsNaN_8U_23U_3_nor_4_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7325" *) _02078_;
  assign IsNaN_8U_23U_3_nor_6_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7326" *) _02079_;
  assign IsNaN_8U_23U_3_nor_8_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7331" *) _02080_;
  assign IsNaN_8U_23U_3_nor_10_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7336" *) _02081_;
  assign _00068_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7354" *) cfg_lut_le_start_rsci_d[22:0];
  assign _02465_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7375" *) reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm;
  assign _02466_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7376" *) reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm;
  assign _02467_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7381" *) FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5;
  assign _02468_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7387" *) reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm;
  assign _02469_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7388" *) reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm;
  assign _02470_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7393" *) FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5;
  assign _02471_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7399" *) reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm;
  assign _02472_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7400" *) reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm;
  assign _02473_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7405" *) FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5;
  assign _02474_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7411" *) reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm;
  assign _02475_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7412" *) reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm;
  assign _02476_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7417" *) FpAdd_8U_23U_2_qr_lpi_1_dfm_5;
  assign IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7456" *) _03746_;
  assign IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7458" *) _03747_;
  assign IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7460" *) _03748_;
  assign IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7462" *) _03749_;
  assign _02477_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7468" *) _01680_;
  assign nor_779_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7472" *) _03752_;
  assign _02478_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7478" *) _01681_;
  assign _02479_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7490" *) _01684_;
  assign _02480_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7498" *) _01685_;
  assign nand_93_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7509" *) _01687_;
  assign _02481_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7511" *) _03756_;
  assign not_tmp_209 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7529" *) _01692_;
  assign not_tmp_222 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7535" *) _01695_;
  assign not_tmp_235 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7539" *) _01697_;
  assign or_tmp_380 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7541" *) _01698_;
  assign not_tmp_248 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7546" *) _01700_;
  assign not_tmp_276 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7561" *) _01703_;
  assign not_tmp_334 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7581" *) _03786_;
  assign _02482_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7584" *) mux_tmp_475;
  assign not_tmp_394 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7584" *) _03787_;
  assign not_tmp_412 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7585" *) _00016_;
  assign not_tmp_418 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7586" *) _03788_;
  assign not_tmp_422 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7587" *) _03789_;
  assign nand_95_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7588" *) and_dcpl_364;
  assign _02483_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7597" *) main_stage_en_1;
  assign _00034_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7600" *) or_tmp_843;
  assign _00035_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7600" *) mux_616_nl;
  assign _02484_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7604" *) _01707_;
  assign nor_647_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7604" *) _03792_;
  assign nor_641_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7613" *) _03793_;
  assign nor_622_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7616" *) _03794_;
  assign _02485_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7633" *) and_tmp_97;
  assign _02486_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *) _01728_;
  assign _02487_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *) _03801_;
  assign nand_tmp_22 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *) _01729_;
  assign _02488_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7652" *) _01739_;
  assign _02489_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7661" *) and_tmp_130;
  assign not_tmp_800 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7667" *) _01750_;
  assign _02490_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7674" *) chn_lut_out_rsci_bawt;
  assign _02491_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7689" *) lut_lookup_1_if_if_else_acc_nl[9];
  assign _02492_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7690" *) _03808_;
  assign _00036_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7695" *) mux_tmp_1130;
  assign _02493_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7696" *) lut_lookup_2_if_if_else_acc_nl[9];
  assign _02494_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7697" *) _03810_;
  assign _00037_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7703" *) mux_tmp_1143;
  assign _02495_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7704" *) lut_lookup_3_if_if_else_acc_nl[9];
  assign _02496_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7705" *) _03812_;
  assign _00038_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7711" *) mux_tmp_1156;
  assign _02497_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7712" *) lut_lookup_4_if_if_else_acc_nl[9];
  assign _02498_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7713" *) _03814_;
  assign _00039_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7719" *) mux_tmp_1169;
  assign _02499_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7722" *) FpAdd_8U_23U_1_is_a_greater_acc_4_nl[8];
  assign _02500_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7723" *) lut_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  assign _02501_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7724" *) lut_lookup_1_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  assign _02502_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7725" *) FpAdd_8U_23U_2_is_a_greater_acc_nl[8];
  assign _02503_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7726" *) lut_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  assign _02504_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7727" *) FpAdd_8U_23U_1_is_a_greater_acc_6_nl[8];
  assign _02505_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7728" *) lut_lookup_2_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  assign _02506_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7729" *) FpAdd_8U_23U_2_is_a_greater_acc_1_nl[8];
  assign _02507_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7730" *) lut_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  assign _02508_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7731" *) FpAdd_8U_23U_1_is_a_greater_acc_8_nl[8];
  assign _02509_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7732" *) lut_lookup_3_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  assign _02510_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7733" *) FpAdd_8U_23U_2_is_a_greater_acc_2_nl[8];
  assign _02511_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7734" *) FpAdd_8U_23U_1_is_a_greater_acc_10_nl[8];
  assign _02512_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7735" *) lut_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  assign _02513_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7736" *) lut_lookup_4_FpAdd_8U_23U_2_is_a_greater_oif_equal_tmp;
  assign _02514_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7737" *) FpAdd_8U_23U_2_is_a_greater_acc_3_nl[8];
  assign _02515_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7742" *) reg_cfg_precision_1_sva_st_12_cse_1[0];
  assign _02516_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7754" *) _01767_;
  assign nor_444_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7754" *) _03823_;
  assign _02517_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7759" *) _01768_;
  assign nor_442_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7759" *) _03824_;
  assign _02518_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7764" *) _01769_;
  assign nor_440_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7764" *) _03825_;
  assign _02519_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7769" *) _01770_;
  assign nor_438_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7769" *) _03826_;
  assign _00069_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7774" *) cfg_lut_lo_start_rsci_d[22:0];
  assign _02520_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7789" *) FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm[7:1];
  assign _02521_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7792" *) FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm[7:1];
  assign _02522_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7795" *) FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm[7:1];
  assign _02523_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7798" *) FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm[7:1];
  assign _02524_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7801" *) FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm[7:1];
  assign _02525_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7804" *) FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm[7:1];
  assign _02526_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7807" *) FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm[7:1];
  assign _02527_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7810" *) FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm[7:1];
  assign _02528_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7814" *) _03827_;
  assign _02529_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7817" *) _03828_;
  assign _02530_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7823" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign _02531_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7836" *) _03834_;
  assign _02532_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7838" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _02533_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7843" *) _03836_;
  assign _02534_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7851" *) _03840_;
  assign nor_823_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7852" *) _03842_;
  assign _02535_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7856" *) _03843_;
  assign nor_820_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7856" *) _03845_;
  assign _02536_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7860" *) _03846_;
  assign nor_817_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7861" *) _03848_;
  assign nor_813_cse = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7864" *) _03849_;
  assign nor_814_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7869" *) _03851_;
  assign _02537_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7886" *) _01773_;
  assign _02538_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7988" *) lut_lookup_le_miss_1_sva;
  assign _02539_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7989" *) lut_lookup_le_miss_2_sva;
  assign _02540_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7990" *) lut_lookup_le_miss_3_sva;
  assign _02541_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7991" *) lut_lookup_le_miss_sva;
  assign _02542_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7992" *) lut_lookup_lo_miss_1_sva;
  assign _02543_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7993" *) lut_lookup_lo_miss_2_sva;
  assign _02544_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7994" *) lut_lookup_lo_miss_3_sva;
  assign _02545_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7995" *) lut_lookup_lo_miss_sva;
  assign _02546_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8087" *) and_dcpl_74;
  assign _02547_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8095" *) main_stage_v_1_mx0c1;
  assign _02548_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8197" *) _03854_;
  assign _02549_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8211" *) _03855_;
  assign _02550_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8217" *) _03856_;
  assign _02551_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8225" *) main_stage_v_2_mx0c1;
  assign _02552_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8310" *) reg_lut_lookup_1_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign _02553_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8363" *) reg_lut_lookup_2_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign _02554_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8412" *) reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign _02555_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8443" *) reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign _02556_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8454" *) main_stage_v_3_mx0c1;
  assign _02557_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8503" *) mux_39_nl;
  assign _02558_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8515" *) mux_1219_nl;
  assign _02559_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8526" *) _03881_;
  assign _02560_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8558" *) mux_1224_nl;
  assign _02561_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8676" *) mux_69_nl;
  assign _02562_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8687" *) mux_82_nl;
  assign _02563_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8724" *) mux_89_nl;
  assign _02564_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8735" *) mux_1226_nl;
  assign _02565_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8746" *) _03884_;
  assign _02566_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8778" *) mux_1230_nl;
  assign _02567_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8835" *) mux_131_nl;
  assign _02568_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8872" *) mux_138_nl;
  assign _02569_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8883" *) mux_1232_nl;
  assign _02570_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8894" *) _03887_;
  assign _02571_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8915" *) _03889_;
  assign _02572_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8927" *) mux_1237_nl;
  assign _02573_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8969" *) mux_167_nl;
  assign _02574_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8992" *) mux_174_nl;
  assign _02575_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9003" *) mux_1239_nl;
  assign _02576_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9014" *) _03893_;
  assign _02577_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9035" *) _03895_;
  assign _02578_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9047" *) mux_1244_nl;
  assign _02579_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9089" *) mux_211_nl;
  assign _02580_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9112" *) main_stage_v_4_mx0c1;
  assign _02581_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9129" *) mux_218_nl;
  assign _02582_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9185" *) lut_lookup_if_else_else_slc_10_mdf_sva_3;
  assign _02583_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9191" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_3;
  assign _02584_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9197" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_3;
  assign _02585_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9215" *) cfg_lut_le_index_select_1_sva_6[0];
  assign _02586_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9235" *) cfg_lut_lo_index_select_1_sva_6[0];
  assign _02587_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9255" *) mux_231_nl;
  assign _02588_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9315" *) mux_244_nl;
  assign _02589_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9375" *) mux_256_nl;
  assign _02590_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9434" *) main_stage_v_5_mx0c1;
  assign _02591_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9491" *) lut_lookup_if_if_lor_5_lpi_1_dfm_4;
  assign _02592_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9494" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_4;
  assign _02593_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9500" *) lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign _02594_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9506" *) lut_lookup_if_if_lor_6_lpi_1_dfm_4;
  assign _02595_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9509" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_4;
  assign _02596_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9515" *) lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign _02597_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9520" *) lut_lookup_if_if_lor_7_lpi_1_dfm_4;
  assign _02598_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9523" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_4;
  assign _02599_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9529" *) lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign _02600_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9534" *) lut_lookup_if_if_lor_1_lpi_1_dfm_4;
  assign _02601_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9537" *) lut_lookup_if_else_else_slc_10_mdf_sva_4;
  assign _02602_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9543" *) lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign _02603_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9617" *) mux_269_nl;
  assign _02604_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9633" *) mux_274_nl;
  assign _02605_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9687" *) mux_281_nl;
  assign _02606_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9763" *) mux_296_nl;
  assign _02607_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9771" *) mux_297_nl;
  assign _02608_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9797" *) mux_301_nl;
  assign _02609_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9805" *) mux_303_nl;
  assign _02610_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9841" *) mux_310_nl;
  assign _02611_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9876" *) mux_320_nl;
  assign _02612_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9885" *) mux_322_nl;
  assign _02613_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9893" *) mux_325_nl;
  assign _02614_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9939" *) mux_334_nl;
  assign _02615_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9964" *) mux_344_nl;
  assign _02616_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9973" *) mux_346_nl;
  assign _02617_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9981" *) mux_349_nl;
  assign _02618_ = and_551_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10307" *) lut_lookup_or_17_rgt;
  assign _02619_ = _02618_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10307" *) lut_lookup_or_18_rgt;
  assign _02620_ = and_559_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10318" *) lut_lookup_and_126_rgt;
  assign _02621_ = _02620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10319" *) lut_lookup_and_127_rgt;
  assign _02622_ = _02621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10319" *) and_564_rgt;
  assign _02623_ = and_566_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10329" *) lut_lookup_and_124_rgt;
  assign _02624_ = _02623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10329" *) lut_lookup_and_125_rgt;
  assign _02625_ = and_570_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10340" *) lut_lookup_and_122_rgt;
  assign _02626_ = _02625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10341" *) lut_lookup_and_123_rgt;
  assign _02627_ = _02626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10341" *) and_564_rgt;
  assign _02628_ = and_576_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10351" *) lut_lookup_and_120_rgt;
  assign _02629_ = _02628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10351" *) lut_lookup_and_121_rgt;
  assign _02630_ = and_580_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10362" *) lut_lookup_and_118_rgt;
  assign _02631_ = _02630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10363" *) lut_lookup_and_119_rgt;
  assign _02632_ = _02631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10363" *) and_586_rgt;
  assign _02633_ = and_588_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10373" *) lut_lookup_or_rgt;
  assign _02634_ = _02633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10373" *) lut_lookup_or_16_rgt;
  assign _02635_ = and_595_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10384" *) lut_lookup_and_112_rgt;
  assign _02636_ = _02635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10385" *) lut_lookup_and_113_rgt;
  assign _02637_ = _02636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10385" *) and_586_rgt;
  assign _02638_ = nor_874_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10673" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _02639_ = and_896_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10744" *) cfg_lut_le_function_1_sva_st_41;
  assign _02640_ = _02639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10744" *) _02115_;
  assign _02641_ = _00985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10789" *) and_653_rgt;
  assign _02642_ = _02639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10892" *) _02121_;
  assign _02643_ = _01011_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10921" *) and_661_rgt;
  assign _02644_ = _02639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11012" *) _02127_;
  assign _02645_ = _01037_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11029" *) and_668_rgt;
  assign _02646_ = _02639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11138" *) _02132_;
  assign _02647_ = _01064_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11155" *) and_676_rgt;
  assign _02648_ = and_427_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11218" *) and_679_rgt;
  assign or_2081_nl = nor_874_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12026" *) or_tmp_1663;
  assign _02649_ = _00001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12028" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
  assign or_1931_nl = _02649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12028" *) _02168_;
  assign _02650_ = nor_792_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12030" *) cfg_lut_le_function_1_sva_st_41;
  assign _02651_ = _02650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12031" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _02652_ = _02651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12031" *) _02169_;
  assign FpAdd_8U_23U_o_expo_or_3_nl = FpAdd_8U_23U_and_51_ssc | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12038" *) _02170_;
  assign or_1941_nl = reg_cfg_precision_1_sva_st_13_cse_1[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12040" *) _02171_;
  assign or_829_nl = IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12050" *) IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
  assign _02653_ = or_829_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12050" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5;
  assign _02654_ = _02653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12050" *) or_tmp_101;
  assign _02655_ = IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12052" *) FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5;
  assign _02656_ = _02655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12052" *) IsNaN_8U_23U_8_land_2_lpi_1_dfm_7;
  assign _02657_ = _02656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12052" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_7;
  assign _02658_ = _02657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12053" *) _00001_;
  assign _02659_ = _02658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12053" *) or_1857_cse;
  assign _02660_ = IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12055" *) nor_13_cse;
  assign _02661_ = _02660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12056" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5;
  assign _02662_ = _02661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12056" *) IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
  assign _02663_ = _02662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12056" *) _00000_;
  assign _02664_ = IsNaN_8U_23U_7_land_1_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12060" *) IsNaN_8U_23U_8_land_2_lpi_1_dfm_7;
  assign _02665_ = _02664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12060" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_6;
  assign _02666_ = _02665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12060" *) FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5;
  assign or_114_nl = or_829_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12075" *) or_tmp_101;
  assign _02667_ = FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12078" *) IsNaN_8U_23U_8_land_2_lpi_1_dfm_7;
  assign _02668_ = _02667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12078" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_7;
  assign _02669_ = _02668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12078" *) _00001_;
  assign or_118_nl = _02669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12078" *) or_1857_cse;
  assign or_120_nl = or_66_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12082" *) IsNaN_8U_23U_7_land_lpi_1_dfm_6;
  assign or_125_nl = or_1857_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12085" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_7;
  assign or_40_nl = _02173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12091" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign or_2080_nl = nor_874_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12096" *) or_tmp_1674;
  assign _02670_ = _00001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12098" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_3;
  assign or_1948_nl = _02670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12098" *) _02174_;
  assign _02671_ = _02650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12101" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  assign _02672_ = _02671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12101" *) _02175_;
  assign FpAdd_8U_23U_o_expo_or_2_nl = FpAdd_8U_23U_and_53_ssc | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12107" *) _02176_;
  assign _02673_ = lut_lookup_2_FpMantRNE_49U_24U_else_and_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12108" *) nor_855_cse;
  assign _02674_ = nor_31_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12116" *) _00000_;
  assign _02675_ = _02674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12117" *) or_66_cse;
  assign _02676_ = _02675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12117" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5;
  assign _02677_ = _02676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12118" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_6;
  assign _02678_ = _02677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12118" *) IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
  assign or_tmp_63 = _00001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12119" *) or_1857_cse;
  assign _02679_ = or_tmp_63 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12120" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_7;
  assign _02680_ = _02679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12120" *) IsNaN_8U_23U_8_land_2_lpi_1_dfm_7;
  assign _02681_ = _02680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12121" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_6;
  assign _02682_ = _02681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12121" *) FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5;
  assign _02683_ = IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12123" *) nor_31_cse;
  assign _02684_ = _02683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12124" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5;
  assign _02685_ = _02684_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12124" *) IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
  assign _02686_ = _02685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12124" *) _00000_;
  assign _02687_ = IsNaN_8U_23U_7_land_2_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12128" *) IsNaN_8U_23U_8_land_2_lpi_1_dfm_7;
  assign _02688_ = _02687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12128" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_6;
  assign _02689_ = _02688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12128" *) FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5;
  assign _02690_ = _02687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12144" *) FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5;
  assign or_184_nl = _02178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12144" *) lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign or_2079_nl = nor_874_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12155" *) or_tmp_1684;
  assign _02691_ = _00001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12157" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_3;
  assign or_1964_nl = _02691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12157" *) _02179_;
  assign _02692_ = _02650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12160" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  assign _02693_ = _02692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12160" *) _02180_;
  assign FpAdd_8U_23U_o_expo_or_1_nl = FpAdd_8U_23U_and_55_ssc | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12168" *) _02176_;
  assign or_1976_nl = reg_cfg_precision_1_sva_st_13_cse_1[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12170" *) _02181_;
  assign _02694_ = IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12179" *) nor_42_cse;
  assign _02695_ = _02694_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12180" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_6;
  assign _02696_ = _02695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12180" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5;
  assign _02697_ = _02696_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12180" *) _00000_;
  assign _02698_ = _02697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12180" *) or_66_cse;
  assign _02699_ = IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12182" *) FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5;
  assign _02700_ = _02699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12182" *) IsNaN_8U_23U_8_land_3_lpi_1_dfm_5;
  assign _02701_ = _02700_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12182" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_7;
  assign _02702_ = _02701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12183" *) or_1857_cse;
  assign _02703_ = _02702_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12183" *) _00001_;
  assign _02704_ = IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12185" *) nor_42_cse;
  assign _02705_ = _02704_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12186" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5;
  assign _02706_ = _02705_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12186" *) IsNaN_8U_23U_8_land_3_lpi_1_dfm_4;
  assign _02707_ = _02706_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12186" *) _00000_;
  assign _02708_ = IsNaN_8U_23U_7_land_3_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12190" *) IsNaN_8U_23U_8_land_3_lpi_1_dfm_5;
  assign _02709_ = _02708_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12190" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_6;
  assign _02710_ = _02709_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12190" *) FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5;
  assign _02711_ = _02695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12205" *) _00000_;
  assign or_247_nl = _02711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12205" *) or_66_cse;
  assign _02712_ = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12208" *) IsNaN_8U_23U_8_land_3_lpi_1_dfm_5;
  assign _02713_ = _02712_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12208" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_7;
  assign _02714_ = _02713_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12208" *) or_1857_cse;
  assign or_251_nl = _02714_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12209" *) _00001_;
  assign or_2078_nl = nor_874_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12220" *) or_tmp_1697;
  assign _02715_ = _00001_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12222" *) lut_lookup_if_else_else_slc_10_mdf_sva_3;
  assign or_1983_nl = _02715_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12222" *) _02183_;
  assign _02716_ = _02650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12225" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign _02717_ = _02716_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12225" *) _02184_;
  assign FpAdd_8U_23U_o_expo_or_nl = FpAdd_8U_23U_and_57_ssc | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12233" *) _02176_;
  assign or_1995_nl = reg_cfg_precision_1_sva_st_13_cse_1[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12235" *) _02185_;
  assign _02718_ = nor_54_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12244" *) _00000_;
  assign _02719_ = _02718_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12245" *) or_66_cse;
  assign _02720_ = _02719_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12245" *) reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse;
  assign _02721_ = _02720_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12246" *) IsNaN_8U_23U_7_land_lpi_1_dfm_6;
  assign _02722_ = _02721_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12246" *) IsNaN_8U_23U_8_land_lpi_1_dfm_4;
  assign _02723_ = or_tmp_63 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12248" *) IsNaN_8U_23U_7_land_lpi_1_dfm_7;
  assign _02724_ = _02723_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12248" *) IsNaN_8U_23U_8_land_lpi_1_dfm_5;
  assign _02725_ = _02724_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12249" *) IsNaN_8U_23U_7_land_lpi_1_dfm_st_6;
  assign _02726_ = _02725_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12249" *) FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5;
  assign _02727_ = IsNaN_8U_23U_7_land_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12251" *) nor_54_cse;
  assign _02728_ = _02727_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12252" *) reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse;
  assign _02729_ = _02728_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12252" *) IsNaN_8U_23U_8_land_lpi_1_dfm_4;
  assign _02730_ = _02729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12252" *) _00000_;
  assign _02731_ = IsNaN_8U_23U_7_land_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12256" *) IsNaN_8U_23U_8_land_lpi_1_dfm_5;
  assign _02732_ = _02731_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12256" *) IsNaN_8U_23U_7_land_lpi_1_dfm_st_6;
  assign _02733_ = _02732_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12256" *) FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5;
  assign or_856_nl = IsNaN_8U_23U_7_land_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12273" *) IsNaN_8U_23U_8_land_lpi_1_dfm_4;
  assign _02734_ = _02187_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12274" *) lut_lookup_4_FpMantRNE_49U_24U_2_else_and_tmp;
  assign _02735_ = _02188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12274" *) _00000_;
  assign or_306_nl = _02735_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12274" *) or_66_cse;
  assign _02736_ = _02189_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12281" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign or_311_nl = _02736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12281" *) _02190_;
  assign _02737_ = _02191_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12284" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3;
  assign or_315_nl = _02737_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12284" *) not_tmp_209;
  assign _02738_ = cfg_lut_le_function_1_sva_st_41 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12287" *) _02190_;
  assign _02739_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12288" *) not_tmp_209;
  assign _02740_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12290" *) _02190_;
  assign _02741_ = lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12293" *) not_tmp_209;
  assign _02742_ = _02192_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12302" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  assign or_341_nl = _02742_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12302" *) _02193_;
  assign _02743_ = _02194_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12305" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3;
  assign or_346_nl = _02743_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12305" *) not_tmp_222;
  assign _02744_ = cfg_lut_le_function_1_sva_st_41 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12308" *) _02193_;
  assign _02745_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12309" *) not_tmp_222;
  assign _02746_ = IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12311" *) _02193_;
  assign _02747_ = lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12314" *) not_tmp_222;
  assign _02748_ = _02195_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12323" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  assign or_374_nl = _02748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12323" *) _02196_;
  assign _02749_ = cfg_lut_le_function_1_sva_st_41 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12328" *) _02196_;
  assign _02750_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12329" *) not_tmp_235;
  assign _02751_ = IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12331" *) _02196_;
  assign _02752_ = _02197_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12342" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign or_406_nl = _02752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12342" *) _02198_;
  assign _02753_ = _02199_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12345" *) lut_lookup_if_else_else_slc_10_mdf_sva_st_3;
  assign or_411_nl = _02753_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12345" *) not_tmp_248;
  assign _02754_ = cfg_lut_le_function_1_sva_st_41 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12348" *) _02198_;
  assign _02755_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12349" *) not_tmp_248;
  assign _02756_ = IsNaN_8U_23U_1_land_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12351" *) _02198_;
  assign _02757_ = lut_lookup_if_else_else_slc_10_mdf_sva_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12354" *) not_tmp_248;
  assign _02758_ = _02200_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12375" *) lut_lookup_else_if_lor_5_lpi_1_dfm_5;
  assign _02759_ = _02758_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12376" *) _02201_;
  assign _02760_ = _02759_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12376" *) IsNaN_8U_23U_6_land_1_lpi_1_dfm_6;
  assign _02761_ = _02760_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12377" *) lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02762_ = _02761_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12377" *) _00032_;
  assign _02763_ = _02762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12377" *) or_tmp_314;
  assign _02764_ = IsNaN_8U_23U_6_land_1_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12379" *) _02202_;
  assign _02765_ = _02764_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12379" *) lut_lookup_else_if_lor_5_lpi_1_dfm_6;
  assign _02766_ = _02765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12380" *) lut_lookup_else_if_lor_5_lpi_1_dfm_st_3;
  assign _02767_ = _02766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12380" *) _02056_;
  assign _02768_ = _02767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12380" *) _02203_;
  assign _02769_ = lut_lookup_else_if_lor_5_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12383" *) _02201_;
  assign _02770_ = _02769_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12384" *) lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02771_ = _02770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12384" *) _00032_;
  assign _02772_ = _02771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12384" *) or_tmp_314;
  assign _02773_ = lut_lookup_else_if_lor_5_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12386" *) lut_lookup_else_if_lor_5_lpi_1_dfm_st_3;
  assign _02774_ = _02773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12386" *) _02056_;
  assign _02775_ = _02774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12386" *) _02203_;
  assign _02776_ = and_854_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12388" *) _02201_;
  assign _02777_ = _02776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12389" *) lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02778_ = _02777_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12389" *) _00032_;
  assign or_445_nl = _02778_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12389" *) or_tmp_314;
  assign _02779_ = _02776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12392" *) IsNaN_8U_23U_6_land_1_lpi_1_dfm_6;
  assign _02780_ = _02779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12393" *) lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02781_ = _02780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12393" *) _00032_;
  assign _02782_ = _02781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12393" *) or_tmp_314;
  assign _02783_ = IsNaN_8U_23U_6_land_1_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12394" *) or_tmp_447;
  assign _02784_ = _02204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12401" *) IsNaN_8U_23U_10_land_1_lpi_1_dfm_5;
  assign _02785_ = _02784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12401" *) lut_lookup_if_1_lor_5_lpi_1_dfm_4;
  assign _02786_ = _02785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12402" *) _00032_;
  assign _02787_ = _02786_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12402" *) or_tmp_314;
  assign _02788_ = _02205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12404" *) lut_lookup_if_1_lor_5_lpi_1_dfm_5;
  assign _02789_ = _02788_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12404" *) IsNaN_8U_23U_10_land_1_lpi_1_dfm_6;
  assign _02790_ = _02789_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12405" *) lut_lookup_if_1_lor_5_lpi_1_dfm_st_4;
  assign _02791_ = _02790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12406" *) _02057_;
  assign _02792_ = _02791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12406" *) _00010_;
  assign _02793_ = lut_lookup_if_1_lor_5_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12409" *) lut_lookup_if_1_lor_5_lpi_1_dfm_st_4;
  assign _02794_ = _02793_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12409" *) _02057_;
  assign _02795_ = _02794_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12409" *) _00010_;
  assign _02796_ = and_846_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12411" *) lut_lookup_if_1_lor_5_lpi_1_dfm_st_4;
  assign _02797_ = _02796_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12412" *) _02057_;
  assign _02798_ = _02797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12412" *) _00010_;
  assign _02799_ = and_846_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12414" *) IsNaN_8U_23U_10_land_1_lpi_1_dfm_6;
  assign _02800_ = _02799_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12415" *) lut_lookup_if_1_lor_5_lpi_1_dfm_st_4;
  assign _02801_ = _02800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12415" *) _02057_;
  assign or_475_nl = _02801_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12415" *) _00010_;
  assign _02802_ = _02206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12422" *) _02201_;
  assign _02803_ = _02802_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12422" *) IsNaN_8U_23U_6_land_2_lpi_1_dfm_6;
  assign _02804_ = _02803_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12424" *) lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02805_ = _02804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12424" *) lut_lookup_else_if_lor_6_lpi_1_dfm_5;
  assign _02806_ = _02805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12424" *) _00032_;
  assign _02807_ = _02806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12424" *) or_tmp_314;
  assign _02808_ = IsNaN_8U_23U_6_land_2_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12426" *) _02207_;
  assign _02809_ = _02808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12426" *) lut_lookup_else_if_lor_6_lpi_1_dfm_6;
  assign _02810_ = _02809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12427" *) lut_lookup_else_if_lor_6_lpi_1_dfm_st_3;
  assign _02811_ = _02810_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12427" *) cfg_precision_1_sva_st_72[0];
  assign _02812_ = _02811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12427" *) not_tmp_276;
  assign _02813_ = _02201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12430" *) lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02814_ = _02813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12430" *) lut_lookup_else_if_lor_6_lpi_1_dfm_5;
  assign _02815_ = _02814_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12430" *) _00032_;
  assign _02816_ = _02815_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12430" *) or_tmp_314;
  assign _02817_ = lut_lookup_else_if_lor_6_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12432" *) lut_lookup_else_if_lor_6_lpi_1_dfm_st_3;
  assign _02818_ = _02817_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12432" *) cfg_precision_1_sva_st_72[0];
  assign _02819_ = _02818_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12432" *) not_tmp_276;
  assign _02820_ = _00032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12435" *) _02201_;
  assign _02821_ = _02820_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12435" *) or_tmp_314;
  assign _02822_ = _02821_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12436" *) lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02823_ = _02822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12436" *) and_82_cse;
  assign or_1851_cse = _02208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12438" *) lut_lookup_else_unequal_tmp_13;
  assign _02824_ = or_1851_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12438" *) _00010_;
  assign _02825_ = _02824_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12438" *) _02056_;
  assign _02826_ = _02825_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12438" *) lut_lookup_else_if_lor_6_lpi_1_dfm_st_3;
  assign _02827_ = _00010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12439" *) _02208_;
  assign _02828_ = _02827_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12440" *) _02056_;
  assign _02829_ = _02828_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12440" *) lut_lookup_else_if_lor_6_lpi_1_dfm_st_3;
  assign _02830_ = _02822_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12445" *) IsNaN_8U_23U_6_land_2_lpi_1_dfm_6;
  assign _02831_ = _02830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12445" *) and_82_cse;
  assign _02832_ = _02826_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12448" *) IsNaN_8U_23U_6_land_2_lpi_1_dfm_7;
  assign _02833_ = _02829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12450" *) IsNaN_8U_23U_6_land_2_lpi_1_dfm_7;
  assign _02834_ = _02209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12458" *) IsNaN_8U_23U_10_land_2_lpi_1_dfm_5;
  assign _02835_ = _02834_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12458" *) lut_lookup_if_1_lor_6_lpi_1_dfm_4;
  assign _02836_ = _02835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12459" *) _00032_;
  assign _02837_ = _02836_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12459" *) or_tmp_314;
  assign _02838_ = IsNaN_8U_23U_10_land_2_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12461" *) _02210_;
  assign _02839_ = _02838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12461" *) lut_lookup_if_1_lor_6_lpi_1_dfm_5;
  assign _02840_ = _02839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12462" *) lut_lookup_if_1_lor_6_lpi_1_dfm_st_4;
  assign _02841_ = _02840_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12462" *) _02057_;
  assign _02842_ = _02841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12462" *) _00010_;
  assign _02843_ = lut_lookup_if_1_lor_6_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12464" *) _00032_;
  assign or_365_cse = _02843_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12465" *) or_tmp_314;
  assign _02844_ = lut_lookup_if_1_lor_6_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12467" *) lut_lookup_if_1_lor_6_lpi_1_dfm_st_4;
  assign _02845_ = _02844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12467" *) _02057_;
  assign _02846_ = _02845_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12467" *) _00010_;
  assign or_528_nl = IsNaN_8U_23U_10_land_2_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12470" *) or_tmp_522;
  assign _02847_ = _02211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12477" *) lut_lookup_else_if_lor_7_lpi_1_dfm_5;
  assign _02848_ = _02847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12478" *) _02201_;
  assign _02849_ = _02848_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12478" *) IsNaN_8U_23U_6_land_3_lpi_1_dfm_6;
  assign _02850_ = _02849_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12479" *) lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02851_ = _02850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12479" *) _00032_;
  assign _02852_ = _02851_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12479" *) or_tmp_314;
  assign _02853_ = IsNaN_8U_23U_6_land_3_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12481" *) _02212_;
  assign _02854_ = _02853_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12481" *) lut_lookup_else_if_lor_7_lpi_1_dfm_6;
  assign _02855_ = _02854_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12482" *) lut_lookup_else_if_lor_7_lpi_1_dfm_st_3;
  assign _02856_ = _02855_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12482" *) _02056_;
  assign _02857_ = _02856_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12482" *) _02203_;
  assign _02858_ = lut_lookup_else_if_lor_7_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12485" *) _02201_;
  assign _02859_ = _02858_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12486" *) lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02860_ = _02859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12486" *) _00032_;
  assign _02861_ = _02860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12486" *) or_tmp_314;
  assign _02862_ = lut_lookup_else_if_lor_7_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12488" *) lut_lookup_else_if_lor_7_lpi_1_dfm_st_3;
  assign _02863_ = _02862_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12488" *) _02056_;
  assign _02864_ = _02863_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12488" *) _02203_;
  assign _02865_ = and_839_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12490" *) _02201_;
  assign _02866_ = _02865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12491" *) lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02867_ = _02866_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12491" *) _00032_;
  assign or_545_nl = _02867_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12491" *) or_tmp_314;
  assign _02868_ = _02865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12494" *) IsNaN_8U_23U_6_land_3_lpi_1_dfm_6;
  assign _02869_ = _02868_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12495" *) lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02870_ = _02869_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12495" *) _00032_;
  assign _02871_ = _02870_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12495" *) or_tmp_314;
  assign _02872_ = IsNaN_8U_23U_6_land_3_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12496" *) or_tmp_547;
  assign _02873_ = _02213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12499" *) IsNaN_8U_23U_10_land_3_lpi_1_dfm_5;
  assign _02874_ = _02873_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12499" *) lut_lookup_if_1_lor_7_lpi_1_dfm_4;
  assign _02875_ = _02874_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12500" *) _00032_;
  assign _02876_ = _02875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12500" *) or_tmp_314;
  assign _02877_ = _02214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12502" *) lut_lookup_if_1_lor_7_lpi_1_dfm_5;
  assign _02878_ = _02877_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12502" *) IsNaN_8U_23U_10_land_3_lpi_1_dfm_6;
  assign _02879_ = _02878_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12503" *) lut_lookup_if_1_lor_7_lpi_1_dfm_st_4;
  assign _02880_ = _02879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12504" *) _02057_;
  assign _02881_ = _02880_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12504" *) _00010_;
  assign _02882_ = lut_lookup_if_1_lor_7_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12507" *) lut_lookup_if_1_lor_7_lpi_1_dfm_st_4;
  assign _02883_ = _02882_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12507" *) _02057_;
  assign or_566_nl = _02883_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12507" *) _00010_;
  assign _02884_ = and_850_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12509" *) lut_lookup_if_1_lor_7_lpi_1_dfm_st_4;
  assign _02885_ = _02884_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12510" *) _02057_;
  assign or_569_nl = _02885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12510" *) _00010_;
  assign _02886_ = and_850_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12512" *) IsNaN_8U_23U_10_land_3_lpi_1_dfm_6;
  assign _02887_ = _02886_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12513" *) lut_lookup_if_1_lor_7_lpi_1_dfm_st_4;
  assign _02888_ = _02887_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12513" *) _02057_;
  assign or_575_nl = _02888_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12513" *) _00010_;
  assign _02889_ = _02215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12520" *) lut_lookup_else_if_lor_1_lpi_1_dfm_5;
  assign _02890_ = _02889_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12521" *) _02201_;
  assign _02891_ = _02890_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12521" *) IsNaN_8U_23U_6_land_lpi_1_dfm_6;
  assign _02892_ = _02891_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12522" *) lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02893_ = _02892_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12522" *) _00032_;
  assign _02894_ = _02893_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12522" *) or_tmp_314;
  assign _02895_ = IsNaN_8U_23U_6_land_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12524" *) _02216_;
  assign _02896_ = _02895_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12524" *) lut_lookup_else_if_lor_1_lpi_1_dfm_6;
  assign _02897_ = _02896_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12525" *) lut_lookup_else_if_lor_1_lpi_1_dfm_st_3;
  assign _02898_ = _02897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12525" *) _02056_;
  assign _02899_ = _02898_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12525" *) _02203_;
  assign _02900_ = lut_lookup_else_if_lor_1_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12528" *) _02201_;
  assign _02901_ = _02900_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12529" *) lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02902_ = _02901_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12529" *) _00032_;
  assign _02903_ = _02902_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12529" *) or_tmp_314;
  assign _02904_ = lut_lookup_else_if_lor_1_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12531" *) lut_lookup_else_if_lor_1_lpi_1_dfm_st_3;
  assign _02905_ = _02904_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12531" *) _02056_;
  assign _02906_ = _02905_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12531" *) _02203_;
  assign _02907_ = and_835_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12533" *) _02201_;
  assign _02908_ = _02907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12534" *) lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02909_ = _02908_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12534" *) _00032_;
  assign or_596_nl = _02909_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12534" *) or_tmp_314;
  assign _02910_ = _02907_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12537" *) IsNaN_8U_23U_6_land_lpi_1_dfm_6;
  assign _02911_ = _02910_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12538" *) lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _02912_ = _02911_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12538" *) _00032_;
  assign _02913_ = _02912_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12538" *) or_tmp_314;
  assign _02914_ = IsNaN_8U_23U_6_land_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12539" *) or_tmp_598;
  assign _02915_ = _02217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12542" *) IsNaN_8U_23U_10_land_lpi_1_dfm_5;
  assign _02916_ = _02915_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12542" *) lut_lookup_if_1_lor_1_lpi_1_dfm_4;
  assign _02917_ = _02916_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12543" *) _00032_;
  assign _02918_ = _02917_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12543" *) or_tmp_314;
  assign _02919_ = _02218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12545" *) lut_lookup_if_1_lor_1_lpi_1_dfm_5;
  assign _02920_ = _02919_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12545" *) IsNaN_8U_23U_10_land_lpi_1_dfm_6;
  assign _02921_ = _02920_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12546" *) lut_lookup_if_1_lor_1_lpi_1_dfm_st_4;
  assign _02922_ = _02921_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12546" *) _02057_;
  assign _02923_ = _02922_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12546" *) _00010_;
  assign _02924_ = lut_lookup_if_1_lor_1_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12549" *) lut_lookup_if_1_lor_1_lpi_1_dfm_st_4;
  assign _02925_ = _02924_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12549" *) _02057_;
  assign or_617_nl = _02925_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12549" *) _00010_;
  assign _02926_ = and_848_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12551" *) lut_lookup_if_1_lor_1_lpi_1_dfm_st_4;
  assign _02927_ = _02926_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12552" *) _02057_;
  assign or_620_nl = _02927_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12552" *) _00010_;
  assign _02928_ = and_848_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12554" *) IsNaN_8U_23U_10_land_lpi_1_dfm_6;
  assign _02929_ = _02928_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12555" *) lut_lookup_if_1_lor_1_lpi_1_dfm_st_4;
  assign _02930_ = _02929_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12555" *) _02057_;
  assign or_625_nl = _02930_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12555" *) _00010_;
  assign _02931_ = lut_lookup_if_else_else_else_asn_mdf_sva_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12560" *) lut_lookup_if_else_else_slc_10_mdf_sva_4;
  assign _02932_ = lut_lookup_4_if_if_else_else_if_acc_nl[3] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12562" *) lut_lookup_4_if_if_else_acc_nl[9];
  assign _02933_ = _02932_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12562" *) lut_lookup_if_if_lor_1_lpi_1_dfm_4;
  assign _02934_ = lut_lookup_if_else_else_else_asn_mdf_2_sva_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12566" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_4;
  assign _02935_ = lut_lookup_2_if_if_else_else_if_acc_nl[3] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12568" *) lut_lookup_2_if_if_else_acc_nl[9];
  assign _02936_ = _02935_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12568" *) lut_lookup_if_if_lor_6_lpi_1_dfm_4;
  assign _02937_ = lut_lookup_if_else_else_else_asn_mdf_1_sva_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12572" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_4;
  assign _02938_ = lut_lookup_1_if_if_else_else_if_acc_nl[3] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12574" *) lut_lookup_1_if_if_else_acc_nl[9];
  assign _02939_ = _02938_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12574" *) lut_lookup_if_if_lor_5_lpi_1_dfm_4;
  assign _02940_ = lut_lookup_if_else_else_else_asn_mdf_3_sva_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12578" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_4;
  assign _02941_ = lut_lookup_3_if_if_else_else_if_acc_nl[3] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12580" *) lut_lookup_3_if_if_else_acc_nl[9];
  assign _02942_ = _02941_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12580" *) lut_lookup_if_if_lor_7_lpi_1_dfm_4;
  assign or_827_nl = main_stage_v_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12612" *) _02227_;
  assign or_186_nl = IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12621" *) IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
  assign _02943_ = nor_193_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12622" *) _02228_;
  assign _02944_ = _02943_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12622" *) _02229_;
  assign or_839_nl = _02944_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12622" *) chn_lut_out_rsci_bawt;
  assign or_850_nl = IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12632" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_6;
  assign or_cse = _02229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12651" *) chn_lut_out_rsci_bawt;
  assign _02945_ = or_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12651" *) _02232_;
  assign _02946_ = IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12692" *) FpAdd_8U_23U_1_mux_61_itm_4;
  assign _02947_ = _02946_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12692" *) IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp;
  assign or_879_nl = _02233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12692" *) or_1857_cse;
  assign _02948_ = lut_lookup_4_if_else_slc_32_svs_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12693" *) nor_792_cse;
  assign _02949_ = _02752_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12695" *) _02184_;
  assign or_880_nl = _02949_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12695" *) lut_lookup_if_else_else_slc_10_mdf_sva_3;
  assign _02950_ = lut_lookup_else_unequal_tmp_12 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12699" *) lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign or_885_nl = _02234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12700" *) or_tmp_314;
  assign or_887_nl = _02235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12702" *) or_tmp_314;
  assign _02951_ = lut_lookup_4_if_else_slc_32_svs_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12704" *) _02236_;
  assign _02952_ = _02237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12706" *) lut_lookup_if_else_else_slc_10_mdf_sva_st_3;
  assign _02953_ = _02952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12706" *) _02238_;
  assign or_888_nl = _02953_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12706" *) lut_lookup_if_else_else_slc_10_mdf_sva_4;
  assign _02954_ = IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12713" *) FpAdd_8U_23U_1_mux_45_itm_4;
  assign _02955_ = _02954_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12713" *) IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp;
  assign or_899_nl = _02239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12713" *) or_1857_cse;
  assign _02956_ = lut_lookup_3_if_else_slc_32_svs_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12714" *) nor_792_cse;
  assign _02957_ = _02748_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12716" *) _02180_;
  assign or_900_nl = _02957_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12716" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_3;
  assign _02958_ = lut_lookup_3_if_else_slc_32_svs_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12722" *) _02236_;
  assign _02959_ = _02240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12724" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3;
  assign _02960_ = _02959_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12724" *) _02241_;
  assign or_907_nl = _02960_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12724" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_4;
  assign _02961_ = IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12730" *) FpAdd_8U_23U_1_mux_29_itm_4;
  assign _02962_ = _02961_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12730" *) IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp;
  assign or_915_nl = _02242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12730" *) or_1857_cse;
  assign _02963_ = lut_lookup_2_if_else_slc_32_svs_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12731" *) nor_792_cse;
  assign _02964_ = _02742_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12733" *) _02175_;
  assign or_916_nl = _02964_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12733" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_3;
  assign _02965_ = lut_lookup_2_if_else_slc_32_svs_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12739" *) _02236_;
  assign _02966_ = _02243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12741" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3;
  assign _02967_ = _02966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12741" *) _02244_;
  assign or_923_nl = _02967_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12741" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_4;
  assign or_931_nl = _02245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12746" *) or_1857_cse;
  assign _02968_ = lut_lookup_1_if_else_slc_32_svs_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12747" *) nor_792_cse;
  assign _02969_ = _02736_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12749" *) _02169_;
  assign or_932_nl = _02969_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12749" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
  assign _02970_ = _02246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12754" *) or_tmp_314;
  assign _02971_ = lut_lookup_1_if_else_slc_32_svs_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12756" *) _02236_;
  assign _02972_ = _02248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12758" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3;
  assign _02973_ = _02972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12758" *) _02249_;
  assign or_939_nl = _02973_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12758" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_4;
  assign _02974_ = FpAdd_8U_23U_2_mux_61_itm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12764" *) and_1138_cse;
  assign _02975_ = _02974_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12764" *) IsZero_8U_23U_8_IsZero_8U_23U_8_nor_3_tmp;
  assign _02976_ = _02250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12765" *) or_1857_cse;
  assign _02977_ = FpAdd_8U_23U_2_mux_45_itm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12768" *) and_1139_cse;
  assign _02978_ = _02977_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12768" *) IsZero_8U_23U_8_IsZero_8U_23U_8_nor_2_tmp;
  assign _02979_ = _02251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12769" *) or_1857_cse;
  assign _02980_ = and_1140_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12773" *) IsZero_8U_23U_8_IsZero_8U_23U_8_nor_1_tmp;
  assign lut_lookup_if_1_lor_6_lpi_1_dfm_mx0w0 = _02980_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12773" *) FpAdd_8U_23U_2_mux_29_itm_3;
  assign _02981_ = lut_lookup_if_1_lor_6_lpi_1_dfm_mx0w0 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12773" *) _00001_;
  assign _02982_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12781" *) _02169_;
  assign _02983_ = _02982_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12781" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
  assign _02984_ = _02983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12782" *) _02252_;
  assign or_990_nl = _02972_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12787" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_4;
  assign _02985_ = IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12801" *) FpAdd_8U_23U_1_mux_13_itm_4;
  assign _02986_ = _02985_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12801" *) mux_1245_nl;
  assign _02987_ = or_932_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12804" *) _02168_;
  assign _02988_ = _02987_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12804" *) cfg_lut_le_function_1_sva_st_41;
  assign _02989_ = _02115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12807" *) cfg_lut_le_function_1_sva_st_41;
  assign _02990_ = _02989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12807" *) _02189_;
  assign _02991_ = _02990_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12808" *) _02168_;
  assign _02992_ = _02991_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12808" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
  assign _02993_ = _02992_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12809" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _02994_ = _02993_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12809" *) _02190_;
  assign _02995_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12811" *) _02253_;
  assign _02996_ = _02995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12812" *) _02254_;
  assign _02997_ = _02996_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12812" *) _02191_;
  assign _02998_ = _02997_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12813" *) _02249_;
  assign _02999_ = _02998_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12813" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3;
  assign _03000_ = _02999_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12814" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_4;
  assign _03001_ = _03000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12815" *) _02255_;
  assign _03002_ = cfg_precision_1_sva_st_71[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12824" *) _02256_;
  assign _03003_ = lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12833" *) lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign or_1045_nl = _03003_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12833" *) _02257_;
  assign _03004_ = nor_792_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12835" *) _02258_;
  assign _03005_ = _03004_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12836" *) FpMantRNE_49U_24U_2_else_carry_1_sva_2;
  assign or_2009_nl = _03005_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12836" *) _02096_;
  assign _03006_ = cfg_precision_1_sva_st_70[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12837" *) _02259_;
  assign or_2007_nl = and_1141_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12839" *) IsZero_8U_23U_8_IsZero_8U_23U_8_nor_tmp;
  assign or_1072_nl = _02966_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12847" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_4;
  assign _03007_ = _02121_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12860" *) cfg_lut_le_function_1_sva_st_41;
  assign _03008_ = _03007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12860" *) _02192_;
  assign _03009_ = _03008_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12861" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_3;
  assign _03010_ = _03009_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12861" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  assign _03011_ = _03010_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12862" *) _02260_;
  assign _03012_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12864" *) _02244_;
  assign _03013_ = _03012_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12864" *) _02194_;
  assign _03014_ = _03013_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12865" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3;
  assign _03015_ = _03014_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12865" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_4;
  assign _03016_ = _03015_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12867" *) _02261_;
  assign _03017_ = cfg_precision_1_sva_st_71[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12873" *) _02262_;
  assign _03018_ = lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12880" *) lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign or_1113_nl = _03018_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12880" *) _02263_;
  assign _03019_ = _02264_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12883" *) FpMantRNE_49U_24U_2_else_carry_2_sva_2;
  assign _03020_ = _03019_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12883" *) _02097_;
  assign or_1142_nl = _02959_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12894" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_4;
  assign _03021_ = _02127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12907" *) cfg_lut_le_function_1_sva_st_41;
  assign _03022_ = _03021_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12907" *) _02195_;
  assign _03023_ = _03022_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12908" *) _02179_;
  assign _03024_ = _03023_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12908" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_3;
  assign _03025_ = _03024_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12909" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  assign _03026_ = _03025_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12909" *) _02196_;
  assign _03027_ = _02265_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12911" *) cfg_lut_le_function_1_sva_st_42;
  assign _03028_ = _03027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12911" *) _02241_;
  assign _03029_ = _03028_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12912" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3;
  assign _03030_ = _03029_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12912" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_4;
  assign _03031_ = _03030_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12914" *) _02266_;
  assign _03032_ = cfg_precision_1_sva_st_71[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12920" *) _02267_;
  assign _03033_ = lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12927" *) lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign or_1183_nl = _03033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12927" *) _02268_;
  assign _03034_ = nor_792_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12929" *) _02269_;
  assign _03035_ = _03034_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12930" *) FpMantRNE_49U_24U_2_else_carry_3_sva_2;
  assign _03036_ = _03035_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12930" *) _02098_;
  assign _03037_ = _02269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12932" *) FpMantRNE_49U_24U_2_else_carry_3_sva_2;
  assign _03038_ = _03037_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12932" *) _02098_;
  assign or_2025_nl = and_1139_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12933" *) IsZero_8U_23U_8_IsZero_8U_23U_8_nor_2_tmp;
  assign _03039_ = cfg_precision_1_sva_st_71[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12939" *) _02270_;
  assign _03040_ = IsNaN_8U_23U_1_land_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12944" *) _02184_;
  assign _03041_ = _03040_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12944" *) lut_lookup_if_else_else_slc_10_mdf_sva_3;
  assign _03042_ = _03041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12945" *) _02271_;
  assign or_1213_nl = _02952_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12950" *) lut_lookup_if_else_else_slc_10_mdf_sva_4;
  assign or_2087_nl = or_1202_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12962" *) cfg_precision_1_sva_st_71[0];
  assign _03043_ = _02132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12967" *) cfg_lut_le_function_1_sva_st_41;
  assign _03044_ = _03043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12967" *) _02197_;
  assign _03045_ = _03044_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12968" *) _02183_;
  assign _03046_ = _03045_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12968" *) lut_lookup_if_else_else_slc_10_mdf_sva_3;
  assign _03047_ = _03046_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12969" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign _03048_ = _03047_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12969" *) _02198_;
  assign _03049_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12971" *) _02238_;
  assign _03050_ = _03049_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12971" *) _02272_;
  assign _03051_ = _03050_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12972" *) _02235_;
  assign _03052_ = _03051_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12972" *) _02199_;
  assign _03053_ = _03052_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12973" *) lut_lookup_if_else_else_slc_10_mdf_sva_4;
  assign _03054_ = _03053_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12973" *) lut_lookup_if_else_else_slc_10_mdf_sva_st_3;
  assign _03055_ = _03054_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12974" *) _02273_;
  assign _03056_ = lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12988" *) lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign or_1252_nl = _03056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12988" *) _02274_;
  assign _03057_ = nor_792_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12990" *) _02275_;
  assign _03058_ = _03057_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12991" *) FpMantRNE_49U_24U_2_else_carry_sva_2;
  assign _03059_ = _03058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12991" *) _02099_;
  assign _03060_ = _02275_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12993" *) FpMantRNE_49U_24U_2_else_carry_sva_2;
  assign _03061_ = _03060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12993" *) _02099_;
  assign or_2035_nl = and_1138_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12994" *) IsZero_8U_23U_8_IsZero_8U_23U_8_nor_3_tmp;
  assign _03062_ = _00000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12998" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _03063_ = _03062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12998" *) lut_lookup_1_if_else_else_acc_nl[10];
  assign _03064_ = _03063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12999" *) _02276_;
  assign _03065_ = nor_792_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13000" *) _00001_;
  assign _03066_ = _03065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13001" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
  assign _03067_ = _03066_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13001" *) _02168_;
  assign _03068_ = cfg_lut_le_function_1_sva_st_41 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13005" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _03069_ = _03068_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13005" *) _02169_;
  assign _03070_ = _03062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13015" *) lut_lookup_2_if_else_else_acc_nl[10];
  assign _03071_ = _03070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13016" *) _02277_;
  assign _03072_ = _03065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13018" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_3;
  assign _03073_ = _03072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13018" *) _02174_;
  assign _03074_ = cfg_lut_le_function_1_sva_st_41 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13022" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  assign _03075_ = _03074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13022" *) _02175_;
  assign _03076_ = _03062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13031" *) lut_lookup_3_if_else_else_acc_nl[10];
  assign _03077_ = _03076_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13032" *) _02278_;
  assign _03078_ = _03065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13034" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_3;
  assign _03079_ = _03078_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13034" *) _02179_;
  assign _03080_ = cfg_lut_le_function_1_sva_st_41 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13038" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  assign _03081_ = _03080_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13038" *) _02180_;
  assign _03082_ = _03062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13047" *) lut_lookup_4_if_else_else_acc_nl[10];
  assign _03083_ = _03082_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13048" *) _02279_;
  assign _03084_ = _03065_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13050" *) lut_lookup_if_else_else_slc_10_mdf_sva_3;
  assign _03085_ = _03084_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13050" *) _02183_;
  assign _03086_ = cfg_lut_le_function_1_sva_st_41 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13054" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign _03087_ = _03086_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13054" *) _02184_;
  assign _03088_ = and_794_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13064" *) and_795_cse;
  assign _03089_ = _03088_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13065" *) or_1495_cse;
  assign _03090_ = _03089_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13065" *) _02280_;
  assign _03091_ = _02281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13067" *) _00033_;
  assign _03092_ = _03091_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13067" *) or_26_cse;
  assign _03093_ = _03092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13067" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _02376_ = IsNaN_8U_23U_4_nor_itm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13069" *) IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2;
  assign _03094_ = _02376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13069" *) _02281_;
  assign _03095_ = _02282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13069" *) _00033_;
  assign _03096_ = _03095_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13070" *) or_26_cse;
  assign _03097_ = _03096_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13070" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _03098_ = and_795_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13073" *) or_1495_cse;
  assign _03099_ = _03098_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13074" *) _02283_;
  assign _03100_ = _03092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13076" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
  assign _03101_ = _01241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13079" *) or_1495_cse;
  assign _03102_ = _03101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13079" *) _02280_;
  assign _03103_ = _01242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13081" *) _00033_;
  assign _03104_ = _03103_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13081" *) or_26_cse;
  assign _03105_ = and_789_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13083" *) and_795_cse;
  assign _03106_ = _03105_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13084" *) or_1495_cse;
  assign _03107_ = _03106_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13084" *) _02280_;
  assign or_1688_cse = _00033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13086" *) or_26_cse;
  assign _03108_ = or_1688_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13086" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
  assign _03109_ = _03108_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13086" *) IsNaN_8U_23U_8_land_2_lpi_1_dfm_5;
  assign _03110_ = and_787_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13088" *) or_tmp_1360;
  assign _03111_ = or_26_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13090" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _03112_ = _03111_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13090" *) IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
  assign _03113_ = _03112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13090" *) _00033_;
  assign _03114_ = and_789_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13092" *) and_787_cse;
  assign _03115_ = _03114_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13093" *) or_1495_cse;
  assign _03116_ = _03115_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13093" *) _02280_;
  assign _03117_ = or_1688_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13095" *) IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
  assign _03118_ = _03117_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13095" *) IsNaN_8U_23U_8_land_2_lpi_1_dfm_5;
  assign _03119_ = and_784_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13097" *) or_tmp_1360;
  assign _03120_ = or_1688_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13099" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _03121_ = _03120_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13099" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  assign _03122_ = and_789_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13101" *) and_784_cse;
  assign _03123_ = _03122_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13102" *) or_1495_cse;
  assign _03124_ = _03123_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13102" *) _02280_;
  assign _03125_ = or_1688_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13104" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  assign _03126_ = _03125_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13104" *) nor_482_cse;
  assign _03127_ = and_794_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13106" *) and_780_cse;
  assign _03128_ = _03127_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13107" *) or_1495_cse;
  assign _03129_ = _03128_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13107" *) _02280_;
  assign _03130_ = _03092_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13109" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _02384_ = IsNaN_8U_23U_4_nor_3_itm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13111" *) IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2;
  assign _03131_ = _02384_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13111" *) _02281_;
  assign _03132_ = _02284_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13111" *) _00033_;
  assign _03133_ = _03132_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13112" *) or_26_cse;
  assign _03134_ = _03133_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13112" *) IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _03135_ = _02285_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13116" *) IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0;
  assign _03136_ = reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13118" *) _00033_;
  assign _03137_ = _03136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13118" *) _02281_;
  assign _03138_ = _03137_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13118" *) or_26_cse;
  assign _03139_ = _01244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13121" *) or_1495_cse;
  assign _03140_ = _03139_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13121" *) _02280_;
  assign _03141_ = _01245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13123" *) _00033_;
  assign _03142_ = _03141_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13123" *) or_26_cse;
  assign _03143_ = and_789_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13125" *) and_780_cse;
  assign _03144_ = _03143_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13126" *) or_1495_cse;
  assign _03145_ = _03144_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13126" *) _02280_;
  assign _03146_ = or_1688_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13128" *) reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse;
  assign _03147_ = _03146_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13128" *) nor_469_cse;
  assign _03148_ = _02286_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13134" *) lut_lookup_1_if_else_else_acc_nl[10];
  assign _03149_ = _03148_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13134" *) _02287_;
  assign _03150_ = _02168_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13139" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
  assign _03151_ = _03150_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13139" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _03152_ = _03151_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13139" *) _02190_;
  assign _03153_ = _02288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13147" *) lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8];
  assign or_1431_nl = _03153_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13147" *) _02289_;
  assign _03154_ = lut_lookup_2_if_else_else_acc_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13153" *) _02290_;
  assign or_1440_nl = lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13164" *) _02291_;
  assign _03155_ = lut_lookup_3_if_else_else_acc_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13170" *) _02292_;
  assign _03156_ = _02293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13180" *) lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8];
  assign or_1450_nl = _03156_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13180" *) _02294_;
  assign _03157_ = _02295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13186" *) lut_lookup_4_if_else_else_acc_nl[10];
  assign _03158_ = _03157_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13186" *) _02296_;
  assign _03159_ = _02183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13190" *) lut_lookup_if_else_else_slc_10_mdf_sva_3;
  assign _03160_ = _03159_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13190" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign _03161_ = _03160_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13190" *) _02198_;
  assign or_1458_nl = lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13199" *) _02297_;
  assign or_1830_nl = reg_cfg_lut_le_function_1_sva_st_20_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13202" *) not_tmp_800;
  assign or_1460_nl = nor_190_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13205" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign _03162_ = reg_cfg_lut_le_function_1_sva_st_19_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13209" *) _02298_;
  assign _03163_ = _00033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13214" *) _02300_;
  assign _03164_ = _03163_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13214" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign _03165_ = _03164_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13214" *) _02301_;
  assign _03166_ = _00033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13219" *) _02302_;
  assign _03167_ = _03166_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13219" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign _03168_ = _03167_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13219" *) _02303_;
  assign _03169_ = reg_cfg_lut_le_function_1_sva_st_20_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13221" *) _02304_;
  assign _03170_ = lut_lookup_else_if_lor_5_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13236" *) lut_lookup_1_else_if_else_if_acc_nl[3];
  assign or_2088_nl = _03170_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13236" *) _02305_;
  assign _03171_ = lut_lookup_else_if_lor_6_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13249" *) lut_lookup_2_else_if_else_if_acc_nl[3];
  assign or_2089_nl = _03171_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13249" *) _02306_;
  assign _03172_ = lut_lookup_else_if_lor_7_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13262" *) lut_lookup_3_else_if_else_if_acc_nl[3];
  assign or_2090_nl = _03172_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13262" *) _02307_;
  assign _03173_ = lut_lookup_else_if_lor_1_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13273" *) lut_lookup_4_else_if_else_if_acc_nl[3];
  assign _03174_ = _03173_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13273" *) _02308_;
  assign _03175_ = _01287_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01301_;
  assign _03176_ = _01288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01302_;
  assign _03177_ = _01289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01303_;
  assign _03178_ = _01290_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01304_;
  assign _03179_ = _01291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01305_;
  assign _03180_ = _01292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01306_;
  assign _03181_ = _01293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01307_;
  assign _03182_ = _01294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01308_;
  assign _03183_ = _01295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01309_;
  assign _03184_ = _01296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01310_;
  assign _03185_ = _01297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01311_;
  assign _03186_ = _01298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01312_;
  assign _03187_ = _01299_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01313_;
  assign _03188_ = _01300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13289" *) _01314_;
  assign _03189_ = _03175_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01315_;
  assign _03190_ = _03176_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01316_;
  assign _03191_ = _03177_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01317_;
  assign _03192_ = _03178_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01318_;
  assign _03193_ = _03179_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01319_;
  assign _03194_ = _03180_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01320_;
  assign _03195_ = _03181_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01321_;
  assign _03196_ = _03182_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01322_;
  assign _03197_ = _03183_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01323_;
  assign _03198_ = _03184_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01323_;
  assign _03199_ = _03185_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01324_;
  assign _03200_ = _03186_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01325_;
  assign _03201_ = _03187_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01326_;
  assign _03202_ = _03188_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13290" *) _01327_;
  assign _03203_ = _01328_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) _01336_;
  assign _03204_ = _01329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) _01337_;
  assign _03205_ = _01330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) _01338_;
  assign _03206_ = _01331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) _01339_;
  assign _03207_ = _01332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) _01340_;
  assign _03208_ = _01333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) _01341_;
  assign _03209_ = _01334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) _01342_;
  assign _03210_ = _01335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13303" *) _01343_;
  assign _03211_ = _03203_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) _01344_;
  assign _03212_ = _03204_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) _01345_;
  assign _03213_ = _03205_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) _01346_;
  assign _03214_ = _03206_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) _01347_;
  assign _03215_ = _03207_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) _01348_;
  assign _03216_ = _03208_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) _01349_;
  assign _03217_ = _03209_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) _01350_;
  assign _03218_ = _03210_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13304" *) _01351_;
  assign _03219_ = _03211_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) _01352_;
  assign _03220_ = _03212_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) _01353_;
  assign _03221_ = _03213_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) _01354_;
  assign _03222_ = _03214_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) _01355_;
  assign _03223_ = _03215_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) _01356_;
  assign _03224_ = _03216_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) _01357_;
  assign _03225_ = _03217_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) _01358_;
  assign _03226_ = _03218_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13305" *) _01359_;
  assign _03227_ = _01360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *) _01364_;
  assign _03228_ = _01361_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *) _01365_;
  assign _03229_ = _01362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *) _01366_;
  assign _03230_ = _01363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13319" *) _01367_;
  assign _03231_ = _03227_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *) _01368_;
  assign _03232_ = _03228_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *) _01369_;
  assign _03233_ = _03229_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *) _01370_;
  assign _03234_ = _03230_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13320" *) _01371_;
  assign _03235_ = _03231_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *) _01372_;
  assign _03236_ = _03232_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *) _01373_;
  assign _03237_ = _03233_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *) _01374_;
  assign _03238_ = _03234_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13321" *) _01375_;
  assign lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_7_nl = _03235_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *) _01376_;
  assign lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_6_nl = _03236_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *) _01377_;
  assign lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_5_nl = _03237_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *) _01378_;
  assign lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_4_nl = _03238_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13322" *) _01379_;
  assign _03239_ = _01380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *) _01384_;
  assign _03240_ = _01381_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *) _01385_;
  assign _03241_ = _01382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *) _01386_;
  assign _03242_ = _01383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13337" *) _01387_;
  assign _03243_ = _03239_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *) _01388_;
  assign _03244_ = _03240_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *) _01389_;
  assign _03245_ = _03241_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *) _01390_;
  assign _03246_ = _03242_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13338" *) _01391_;
  assign _03247_ = _03243_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *) _01392_;
  assign _03248_ = _03244_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *) _01393_;
  assign _03249_ = _03245_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *) _01394_;
  assign _03250_ = _03246_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13339" *) _01395_;
  assign _03251_ = _03247_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *) _01396_;
  assign _03252_ = _03248_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *) _01397_;
  assign _03253_ = _03249_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *) _01398_;
  assign _03254_ = _03250_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13340" *) _01399_;
  assign _03255_ = _03251_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *) _01400_;
  assign _03256_ = _03252_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *) _01401_;
  assign _03257_ = _03253_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *) _01402_;
  assign _03258_ = _03254_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13341" *) _01403_;
  assign _03259_ = _01404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *) _01408_;
  assign _03260_ = _01405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *) _01409_;
  assign _03261_ = _01406_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *) _01410_;
  assign _03262_ = _01407_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13353" *) _01411_;
  assign _03263_ = _03259_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *) _01412_;
  assign _03264_ = _03260_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *) _01413_;
  assign _03265_ = _03261_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *) _01414_;
  assign _03266_ = _03262_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13354" *) _01415_;
  assign _03267_ = _01416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *) _01420_;
  assign _03268_ = _01417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *) _01421_;
  assign _03269_ = _01418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *) _01422_;
  assign _03270_ = _01419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13367" *) _01423_;
  assign _03271_ = _03267_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *) _01424_;
  assign _03272_ = _03268_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *) _01425_;
  assign _03273_ = _03269_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *) _01426_;
  assign _03274_ = _03270_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13368" *) _01427_;
  assign _03275_ = _03271_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *) _01428_;
  assign _03276_ = _03272_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *) _01429_;
  assign _03277_ = _03273_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *) _01430_;
  assign _03278_ = _03274_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13369" *) _01431_;
  assign _03279_ = _01432_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *) _01436_;
  assign _03280_ = _01433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *) _01437_;
  assign _03281_ = _01434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *) _01438_;
  assign _03282_ = _01435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13381" *) _01439_;
  assign _03283_ = _03279_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *) _01440_;
  assign _03284_ = _03280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *) _01441_;
  assign _03285_ = _03281_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *) _01442_;
  assign _03286_ = _03282_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13382" *) _01443_;
  assign _03287_ = _01444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *) _01448_;
  assign _03288_ = _01445_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *) _01449_;
  assign _03289_ = _01446_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *) _01450_;
  assign _03290_ = _01447_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13397" *) _01451_;
  assign _03291_ = _03287_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *) _01452_;
  assign _03292_ = _03288_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *) _01453_;
  assign _03293_ = _03289_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *) _01454_;
  assign _03294_ = _03290_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13398" *) _01455_;
  assign _03295_ = _03291_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *) _01456_;
  assign _03296_ = _03292_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *) _01457_;
  assign _03297_ = _03293_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *) _01458_;
  assign _03298_ = _03294_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13399" *) _01459_;
  assign _03299_ = _03295_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *) _01460_;
  assign _03300_ = _03296_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *) _01461_;
  assign _03301_ = _03297_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *) _01462_;
  assign _03302_ = _03298_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13400" *) _01463_;
  assign _03303_ = _03299_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *) _01464_;
  assign _03304_ = _03300_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *) _01465_;
  assign _03305_ = _03301_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *) _01466_;
  assign _03306_ = _03302_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13401" *) _01467_;
  assign _03307_ = _01468_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *) _01472_;
  assign _03308_ = _01469_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *) _01473_;
  assign _03309_ = _01470_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *) _01474_;
  assign _03310_ = _01471_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13413" *) _01475_;
  assign _03311_ = _03307_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *) _01476_;
  assign _03312_ = _03308_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *) _01477_;
  assign _03313_ = _03309_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *) _01478_;
  assign _03314_ = _03310_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13414" *) _01479_;
  assign _03315_ = _01480_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) _01488_;
  assign _03316_ = _01481_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) _01489_;
  assign _03317_ = _01482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) _01490_;
  assign _03318_ = _01483_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) _01491_;
  assign _03319_ = _01484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) _01492_;
  assign _03320_ = _01485_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) _01493_;
  assign _03321_ = _01486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) _01494_;
  assign _03322_ = _01487_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13428" *) _01495_;
  assign _03323_ = _03315_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) _01496_;
  assign _03324_ = _03316_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) _01497_;
  assign _03325_ = _03317_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) _01498_;
  assign _03326_ = _03318_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) _01499_;
  assign _03327_ = _03319_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) _01500_;
  assign _03328_ = _03320_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) _01501_;
  assign _03329_ = _03321_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) _01502_;
  assign _03330_ = _03322_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13429" *) _01503_;
  assign _03331_ = _03323_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) _01504_;
  assign _03332_ = _03324_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) _01505_;
  assign _03333_ = _03325_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) _01506_;
  assign _03334_ = _03326_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) _01507_;
  assign _03335_ = _03327_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) _01508_;
  assign _03336_ = _03328_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) _01509_;
  assign _03337_ = _03329_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) _01510_;
  assign _03338_ = _03330_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13430" *) _01511_;
  assign FpAdd_8U_23U_FpAdd_8U_23U_mux1h_2_tmp = _03331_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) _01512_;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_2_tmp = _03332_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) _01513_;
  assign FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7 = _03333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) _01514_;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_5_tmp = _03334_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) _01515_;
  assign FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7 = _03335_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) _01516_;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_8_tmp = _03336_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) _01517_;
  assign FpAdd_8U_23U_o_expo_lpi_1_dfm_7 = _03337_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) _01518_;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_mux1h_11_tmp = _03338_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13431" *) _01519_;
  assign _03339_ = _01520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *) _01524_;
  assign _03340_ = _01521_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *) _01525_;
  assign _03341_ = _01522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *) _01526_;
  assign _03342_ = _01523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13445" *) _01527_;
  assign _03343_ = _03339_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13446" *) _01528_;
  assign _03344_ = _03340_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13446" *) _01528_;
  assign _03345_ = _03341_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13446" *) _01528_;
  assign _03346_ = _03342_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13446" *) _01528_;
  assign _03347_ = _03343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *) _01529_;
  assign _03348_ = _03344_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *) _01530_;
  assign _03349_ = _03345_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *) _01531_;
  assign _03350_ = _03346_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13447" *) _01532_;
  assign lut_lookup_else_else_else_else_mux1h_rgt = _03347_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13448" *) _01533_;
  assign lut_lookup_else_else_else_else_mux1h_1_rgt = _03348_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13448" *) _01533_;
  assign lut_lookup_else_else_else_else_mux1h_2_rgt = _03349_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13448" *) _01533_;
  assign lut_lookup_else_else_else_else_mux1h_3_rgt = _03350_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13448" *) _01533_;
  assign _03351_ = and_dcpl_54 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5452" *) _00010_;
  assign _03352_ = _01534_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5454" *) and_dcpl_59;
  assign _03353_ = _01535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5456" *) and_dcpl_63;
  assign _03354_ = _01536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5458" *) and_dcpl_67;
  assign _03355_ = _01537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5460" *) and_dcpl_71;
  assign _03356_ = or_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5475" *) nor_193_cse;
  assign _03357_ = nor_874_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5496" *) reg_cfg_precision_1_sva_st_12_cse_1[0];
  assign IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_5_cse = _01538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5498" *) and_524_rgt;
  assign _03358_ = reg_cfg_lut_le_function_1_sva_st_19_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5503" *) reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign _03359_ = reg_cfg_lut_le_function_1_sva_st_19_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5512" *) reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign _03360_ = nor_5_cse_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5532" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5;
  assign _03361_ = _03360_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5533" *) IsNaN_8U_23U_4_land_1_lpi_1_dfm_4;
  assign _03362_ = _03361_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5533" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign _03363_ = _03362_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5533" *) _00000_;
  assign _03364_ = _03363_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5533" *) or_66_cse;
  assign _03365_ = IsNaN_8U_23U_3_land_1_lpi_1_dfm_st_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5535" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _03366_ = _03365_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5535" *) FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6;
  assign _03367_ = _03366_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5535" *) IsNaN_8U_23U_3_land_1_lpi_1_dfm_6;
  assign _03368_ = _03367_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5536" *) _00001_;
  assign _03369_ = _03368_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5536" *) or_1857_cse;
  assign _03370_ = lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5540" *) _02330_;
  assign _03371_ = mux_1220_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5556" *) nor_5_cse_1;
  assign _03372_ = _03371_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5556" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign or_1936_cse = _02333_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5557" *) lut_lookup_1_FpMantRNE_49U_24U_else_and_tmp;
  assign _03373_ = nor_874_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5558" *) reg_cfg_precision_1_sva_st_13_cse_1[0];
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_6_cse = _01544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5559" *) and_dcpl_161;
  assign IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_3_aelse_or_3_cse = and_dcpl_148 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5560" *) and_dcpl_162;
  assign _03374_ = lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5564" *) _02335_;
  assign FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse = and_401_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5566" *) and_dcpl_161;
  assign _03375_ = FpAdd_8U_23U_2_int_mant_p1_1_sva_3[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5568" *) and_dcpl_54;
  assign _03376_ = and_364_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5579" *) and_dcpl_148;
  assign IsNaN_8U_23U_1_aelse_IsNaN_8U_23U_1_aelse_or_8_cse = _03376_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5579" *) and_347_rgt;
  assign _03377_ = nor_27_cse_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5580" *) _00000_;
  assign _03378_ = _03377_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5581" *) or_66_cse;
  assign _03379_ = _03378_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5581" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5;
  assign _03380_ = _03379_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5582" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _03381_ = _03380_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5582" *) IsNaN_8U_23U_4_land_2_lpi_1_dfm_5;
  assign _03382_ = or_tmp_63 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5584" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  assign _03383_ = _03382_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5584" *) IsNaN_8U_23U_3_land_2_lpi_1_dfm_7;
  assign _03384_ = _03383_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5585" *) IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_6;
  assign _03385_ = _03384_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5585" *) FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6;
  assign _03386_ = lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5590" *) _02337_;
  assign _03387_ = mux_1227_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5606" *) nor_27_cse_1;
  assign _03388_ = _03387_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5606" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _03389_ = lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5611" *) _02340_;
  assign _03390_ = FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5613" *) and_dcpl_54;
  assign or_48_cse = _02343_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5620" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _03391_ = nor_38_cse_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5621" *) _00000_;
  assign _03392_ = _03391_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5622" *) or_66_cse;
  assign _03393_ = _03392_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5622" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5;
  assign _03394_ = _03393_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5623" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign _03395_ = _03394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5623" *) IsNaN_8U_23U_4_land_3_lpi_1_dfm_5;
  assign _03396_ = or_tmp_63 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5625" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  assign _03397_ = _03396_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5625" *) IsNaN_8U_23U_3_land_3_lpi_1_dfm_7;
  assign _03398_ = _03397_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5626" *) IsNaN_8U_23U_3_land_3_lpi_1_dfm_st_6;
  assign _03399_ = _03398_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5626" *) FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6;
  assign _03400_ = lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5630" *) _02344_;
  assign _03401_ = lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5644" *) _02347_;
  assign _03402_ = FpAdd_8U_23U_2_int_mant_p1_3_sva_3[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5647" *) and_dcpl_54;
  assign _03403_ = nor_50_cse_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5652" *) _00000_;
  assign _03404_ = _03403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5653" *) or_66_cse;
  assign _03405_ = _03404_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5653" *) reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse;
  assign _03406_ = _03405_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5654" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _03407_ = _03406_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5654" *) IsNaN_8U_23U_4_land_lpi_1_dfm_4;
  assign _03408_ = or_tmp_63 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5656" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign _03409_ = _03408_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5656" *) IsNaN_8U_23U_3_land_lpi_1_dfm_6;
  assign _03410_ = _03409_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5657" *) IsNaN_8U_23U_3_land_lpi_1_dfm_st_6;
  assign _03411_ = _03410_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5657" *) FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6;
  assign _03412_ = lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5661" *) _02349_;
  assign _03413_ = lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5675" *) _02352_;
  assign _03414_ = FpAdd_8U_23U_2_int_mant_p1_sva_3[49] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5677" *) and_dcpl_54;
  assign or_312_cse = _00032_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5684" *) or_tmp_314;
  assign lut_lookup_if_else_else_else_else_if_lut_lookup_if_else_else_else_else_if_or_3_cse = and_427_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5686" *) and_428_rgt;
  assign _03415_ = cfg_lut_le_function_1_sva_st_41 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5687" *) _02354_;
  assign _03416_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5688" *) _02355_;
  assign _03417_ = _02112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5692" *) and_1142_cse;
  assign _03418_ = _03417_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5693" *) FpAdd_8U_23U_1_mux_13_itm_4;
  assign _03419_ = _03418_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5693" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp;
  assign _03420_ = _03419_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5693" *) _00001_;
  assign _03421_ = _03420_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5693" *) or_1857_cse;
  assign _03422_ = _02201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5695" *) lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _03423_ = _03422_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5695" *) _00032_;
  assign _03424_ = _03423_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5695" *) or_tmp_314;
  assign FpAdd_8U_23U_1_lut_lookup_else_else_else_or_3_cse = _01561_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5701" *) and_430_rgt;
  assign _03425_ = lut_lookup_if_1_lor_5_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5702" *) _00032_;
  assign or_332_nl = _03425_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5702" *) or_tmp_314;
  assign _03426_ = _02112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5707" *) IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp;
  assign _03427_ = _03426_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5707" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp;
  assign _03428_ = _03427_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5707" *) FpAdd_8U_23U_1_mux_29_itm_4;
  assign _03429_ = _03428_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5708" *) _00001_;
  assign _03430_ = _03429_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5708" *) or_1857_cse;
  assign _03431_ = _02813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5710" *) _00032_;
  assign _03432_ = _03431_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5710" *) or_tmp_314;
  assign _03433_ = _02112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5720" *) IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp;
  assign _03434_ = _03433_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5720" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp;
  assign _03435_ = _03434_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5720" *) FpAdd_8U_23U_1_mux_45_itm_4;
  assign _03436_ = _03435_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5721" *) _00001_;
  assign _03437_ = _03436_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5721" *) or_1857_cse;
  assign _03438_ = _02201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5723" *) lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _03439_ = _03438_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5723" *) _00032_;
  assign _03440_ = _03439_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5723" *) or_tmp_314;
  assign _03441_ = _02112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5731" *) IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp;
  assign _03442_ = _03441_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5731" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp;
  assign _03443_ = _03442_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5732" *) FpAdd_8U_23U_1_mux_61_itm_4;
  assign _03444_ = _03443_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5732" *) _00001_;
  assign _03445_ = _03444_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5732" *) or_1857_cse;
  assign _03446_ = _02201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5734" *) lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _03447_ = _03446_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5734" *) _00032_;
  assign _03448_ = _03447_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5734" *) or_tmp_314;
  assign or_1853_cse = _02201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5744" *) lut_lookup_else_unequal_tmp_18;
  assign or_492_cse = _02201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5759" *) lut_lookup_else_unequal_tmp_12;
  assign _03449_ = and_dcpl_258 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5776" *) and_dcpl_259;
  assign _03450_ = or_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5780" *) _02365_;
  assign _03451_ = and_dcpl_258 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5786" *) and_465_cse;
  assign lut_lookup_else_else_lut_lookup_else_else_or_3_cse = _03451_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5786" *) and_466_cse;
  assign lut_lookup_FpAdd_8U_23U_1_or_11_cse = _01563_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5799" *) and_dcpl_280;
  assign lut_lookup_FpAdd_8U_23U_2_or_10_cse = _01564_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5803" *) and_dcpl_292;
  assign lut_lookup_FpAdd_8U_23U_2_or_9_cse = _01565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5807" *) and_dcpl_300;
  assign lut_lookup_FpAdd_8U_23U_2_or_8_cse = _01566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5809" *) and_dcpl_308;
  assign FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_cse = _01567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5811" *) FpAdd_8U_23U_1_is_a_greater_acc_4_nl[8];
  assign _03452_ = _01569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5814" *) _01571_;
  assign _03453_ = _03452_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5814" *) and_dcpl_314;
  assign IsZero_8U_23U_1_IsZero_8U_23U_4_or_3_cse = and_dcpl_315 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5815" *) and_dcpl_316;
  assign FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_cse = _01573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5819" *) FpAdd_8U_23U_2_is_a_greater_acc_nl[8];
  assign _03454_ = _01574_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5821" *) and_dcpl_314;
  assign FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_1_cse = _01576_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5823" *) FpAdd_8U_23U_1_is_a_greater_acc_6_nl[8];
  assign FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_1_cse = _01577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5827" *) FpAdd_8U_23U_2_is_a_greater_acc_1_nl[8];
  assign FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_2_cse = _01578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5829" *) FpAdd_8U_23U_1_is_a_greater_acc_8_nl[8];
  assign FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_2_cse = _01579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5831" *) FpAdd_8U_23U_2_is_a_greater_acc_2_nl[8];
  assign FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_3_cse = _01580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5834" *) FpAdd_8U_23U_1_is_a_greater_acc_10_nl[8];
  assign FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_3_cse = _01581_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5836" *) FpAdd_8U_23U_2_is_a_greater_acc_3_nl[8];
  assign _03455_ = _01582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5841" *) and_525_rgt;
  assign _03456_ = and_527_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5845" *) and_529_rgt;
  assign _03457_ = _03456_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5846" *) and_525_rgt;
  assign lut_lookup_or_17_rgt = _01587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5853" *) _01588_;
  assign lut_lookup_or_18_rgt = _01589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5855" *) _01590_;
  assign or_tmp_6 = _02280_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5858" *) or_1495_cse;
  assign or_1689_cse = _00000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5859" *) or_66_cse;
  assign or_849_cse = _00033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5888" *) reg_cfg_precision_1_sva_st_12_cse_1[0];
  assign or_1696_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5890" *) _02281_;
  assign lut_lookup_or_rgt = _01599_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5895" *) _01600_;
  assign lut_lookup_or_16_rgt = _01601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5897" *) _01602_;
  assign _03458_ = and_604_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5905" *) and_606_rgt;
  assign _03459_ = _03458_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5905" *) and_dcpl_403;
  assign IsNaN_8U_23U_5_IsNaN_8U_23U_6_aelse_or_2_cse = _03459_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5905" *) and_dcpl_405;
  assign mux_670_cse = mux_1285_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5908" *) _02112_;
  assign _03460_ = _02389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5912" *) or_tmp_314;
  assign _03461_ = FpAdd_8U_23U_2_mux_13_itm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5926" *) and_1141_cse;
  assign or_969_cse = _03461_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5926" *) IsZero_8U_23U_8_IsZero_8U_23U_8_nor_tmp;
  assign or_978_cse = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5927" *) _00032_;
  assign mux_745_cse = mux_1282_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5930" *) cfg_lut_le_function_1_sva_st_41;
  assign _03462_ = nor_610_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5944" *) _00032_;
  assign _03463_ = _02394_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5964" *) _02059_;
  assign _03464_ = _02112_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5965" *) or_1857_cse;
  assign _03465_ = _02201_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5966" *) or_tmp_314;
  assign _03466_ = lut_lookup_1_if_else_else_else_else_acc_nl[32] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5975" *) cfg_lut_le_function_1_sva_st_41;
  assign _03467_ = _03466_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5975" *) and_896_cse;
  assign _03468_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5977" *) lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _03469_ = _03468_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5977" *) _02236_;
  assign _03470_ = _02989_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5980" *) and_896_cse;
  assign _03471_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5982" *) _02395_;
  assign _03472_ = IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6013" *) _02175_;
  assign _03473_ = _03472_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6013" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_3;
  assign _03474_ = _03473_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6014" *) _02397_;
  assign _03475_ = lut_lookup_2_if_else_else_else_else_acc_nl[32] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6033" *) cfg_lut_le_function_1_sva_st_41;
  assign _03476_ = _03475_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6033" *) and_896_cse;
  assign _03477_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6035" *) lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _03478_ = _03477_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6035" *) _02236_;
  assign _03479_ = _03007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6038" *) and_896_cse;
  assign _03480_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6040" *) _02399_;
  assign _03481_ = IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6059" *) _02180_;
  assign _03482_ = _03481_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6059" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_3;
  assign _03483_ = _03482_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6060" *) _02401_;
  assign _03484_ = lut_lookup_3_if_else_else_else_else_acc_nl[32] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6078" *) cfg_lut_le_function_1_sva_st_41;
  assign _03485_ = _03484_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6078" *) and_896_cse;
  assign _03486_ = lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6080" *) cfg_lut_le_function_1_sva_st_42;
  assign _03487_ = _03486_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6080" *) _02236_;
  assign _03488_ = _03021_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6083" *) and_896_cse;
  assign _03489_ = _02403_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6085" *) cfg_lut_le_function_1_sva_st_42;
  assign _03490_ = _03489_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6085" *) _02236_;
  assign _03491_ = lut_lookup_4_if_else_else_else_else_acc_nl[32] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6120" *) cfg_lut_le_function_1_sva_st_41;
  assign _03492_ = _03491_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6120" *) and_896_cse;
  assign _03493_ = IsNaN_8U_23U_6_land_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6121" *) _02236_;
  assign _03494_ = _03043_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6124" *) and_896_cse;
  assign _03495_ = cfg_lut_le_function_1_sva_st_42 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6125" *) _02272_;
  assign _03496_ = cfg_precision_1_sva_st_71[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6131" *) _00032_;
  assign _02383_ = IsNaN_8U_23U_8_nor_2_itm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6157" *) IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_2;
  assign _03497_ = and_784_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6158" *) _02280_;
  assign _03498_ = _03497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6158" *) or_1495_cse;
  assign _03499_ = _00033_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6160" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  assign _03500_ = _03499_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6160" *) or_26_cse;
  assign _02387_ = IsNaN_8U_23U_8_nor_3_itm_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6164" *) IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_3_itm_2;
  assign _03501_ = or_tmp_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6166" *) IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0;
  assign _03502_ = _03136_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6168" *) or_26_cse;
  assign _03503_ = IsNaN_8U_23U_3_nor_8_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6191" *) _02064_;
  assign _03504_ = IsNaN_8U_23U_3_nor_6_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6192" *) _02065_;
  assign _03505_ = FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6199" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[1];
  assign _03506_ = _03505_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6199" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[2];
  assign _03507_ = _03506_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6200" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[3];
  assign _03508_ = _03507_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6200" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[4];
  assign _03509_ = _03508_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6201" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[5];
  assign _03510_ = _03509_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6201" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[6];
  assign _03511_ = _03510_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6202" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[7];
  assign _03512_ = _03511_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6202" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[8];
  assign _03513_ = _03512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6203" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[9];
  assign _03514_ = _03513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6203" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[10];
  assign _03515_ = _03514_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6204" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[11];
  assign _03516_ = _03515_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6204" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[12];
  assign _03517_ = _03516_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6205" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[13];
  assign _03518_ = _03517_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6205" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[14];
  assign _03519_ = _03518_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6206" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[15];
  assign _03520_ = _03519_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6206" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[16];
  assign _03521_ = _03520_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6207" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[17];
  assign _03522_ = _03521_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6207" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[18];
  assign _03523_ = _03522_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6208" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[19];
  assign _03524_ = _03523_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6208" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[20];
  assign _03525_ = _03524_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6209" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[21];
  assign _03526_ = _03525_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6209" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[22];
  assign _03527_ = _03526_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6210" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[23];
  assign _03528_ = _03527_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6210" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[25];
  assign _03529_ = FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6219" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[1];
  assign _03530_ = _03529_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6219" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[2];
  assign _03531_ = _03530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6220" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[3];
  assign _03532_ = _03531_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6220" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[4];
  assign _03533_ = _03532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6221" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[5];
  assign _03534_ = _03533_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6221" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[6];
  assign _03535_ = _03534_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6222" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[7];
  assign _03536_ = _03535_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6222" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[8];
  assign _03537_ = _03536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6223" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[9];
  assign _03538_ = _03537_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6223" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[10];
  assign _03539_ = _03538_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6224" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[11];
  assign _03540_ = _03539_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6224" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[12];
  assign _03541_ = _03540_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6225" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[13];
  assign _03542_ = _03541_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6225" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[14];
  assign _03543_ = _03542_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6226" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[15];
  assign _03544_ = _03543_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6226" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[16];
  assign _03545_ = _03544_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6227" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[17];
  assign _03546_ = _03545_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6227" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[18];
  assign _03547_ = _03546_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6228" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[19];
  assign _03548_ = _03547_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6228" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[20];
  assign _03549_ = _03548_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6229" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[21];
  assign _03550_ = _03549_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6229" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[22];
  assign _03551_ = _03550_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6230" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[23];
  assign _03552_ = _03551_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6230" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[25];
  assign _03553_ = FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6239" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[1];
  assign _03554_ = _03553_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6239" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[2];
  assign _03555_ = _03554_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6240" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[3];
  assign _03556_ = _03555_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6240" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[4];
  assign _03557_ = _03556_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6241" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[5];
  assign _03558_ = _03557_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6241" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[6];
  assign _03559_ = _03558_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6242" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[7];
  assign _03560_ = _03559_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6242" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[8];
  assign _03561_ = _03560_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6243" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[9];
  assign _03562_ = _03561_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6243" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[10];
  assign _03563_ = _03562_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6244" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[11];
  assign _03564_ = _03563_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6244" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[12];
  assign _03565_ = _03564_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6245" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[13];
  assign _03566_ = _03565_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6245" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[14];
  assign _03567_ = _03566_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6246" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[15];
  assign _03568_ = _03567_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6246" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[16];
  assign _03569_ = _03568_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6247" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[17];
  assign _03570_ = _03569_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6247" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[18];
  assign _03571_ = _03570_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6248" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[19];
  assign _03572_ = _03571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6248" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[20];
  assign _03573_ = _03572_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6249" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[21];
  assign _03574_ = _03573_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6249" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[22];
  assign _03575_ = _03574_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6250" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[23];
  assign _03576_ = _03575_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6250" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[25];
  assign _03577_ = FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6259" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[1];
  assign _03578_ = _03577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6259" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[2];
  assign _03579_ = _03578_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6260" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[3];
  assign _03580_ = _03579_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6260" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[4];
  assign _03581_ = _03580_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6261" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[5];
  assign _03582_ = _03581_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6261" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[6];
  assign _03583_ = _03582_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6262" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[7];
  assign _03584_ = _03583_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6262" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[8];
  assign _03585_ = _03584_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6263" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[9];
  assign _03586_ = _03585_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6263" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[10];
  assign _03587_ = _03586_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6264" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[11];
  assign _03588_ = _03587_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6264" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[12];
  assign _03589_ = _03588_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6265" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[13];
  assign _03590_ = _03589_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6265" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[14];
  assign _03591_ = _03590_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6266" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[15];
  assign _03592_ = _03591_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6266" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[16];
  assign _03593_ = _03592_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6267" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[17];
  assign _03594_ = _03593_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6267" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[18];
  assign _03595_ = _03594_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6268" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[19];
  assign _03596_ = _03595_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6268" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[20];
  assign _03597_ = _03596_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6269" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[21];
  assign _03598_ = _03597_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6269" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[22];
  assign _03599_ = _03598_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6270" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[23];
  assign _03600_ = _03599_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6270" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[25];
  assign _03601_ = FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6279" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[1];
  assign _03602_ = _03601_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6279" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[2];
  assign _03603_ = _03602_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6280" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[3];
  assign _03604_ = _03603_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6280" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[4];
  assign _03605_ = _03604_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6281" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[5];
  assign _03606_ = _03605_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6281" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[6];
  assign _03607_ = _03606_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6282" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[7];
  assign _03608_ = _03607_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6282" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[8];
  assign _03609_ = _03608_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6283" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[9];
  assign _03610_ = _03609_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6283" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[10];
  assign _03611_ = _03610_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6284" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[11];
  assign _03612_ = _03611_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6284" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[12];
  assign _03613_ = _03612_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6285" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[13];
  assign _03614_ = _03613_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6285" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[14];
  assign _03615_ = _03614_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6286" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[15];
  assign _03616_ = _03615_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6286" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[16];
  assign _03617_ = _03616_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6287" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[17];
  assign _03618_ = _03617_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6287" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[18];
  assign _03619_ = _03618_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6288" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[19];
  assign _03620_ = _03619_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6288" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[20];
  assign _03621_ = _03620_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6289" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[21];
  assign _03622_ = _03621_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6289" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[22];
  assign _03623_ = _03622_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6290" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[23];
  assign _03624_ = _03623_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6290" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[25];
  assign _03625_ = FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6299" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[1];
  assign _03626_ = _03625_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6299" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[2];
  assign _03627_ = _03626_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6300" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[3];
  assign _03628_ = _03627_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6300" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[4];
  assign _03629_ = _03628_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6301" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[5];
  assign _03630_ = _03629_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6301" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[6];
  assign _03631_ = _03630_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6302" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[7];
  assign _03632_ = _03631_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6302" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[8];
  assign _03633_ = _03632_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6303" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[9];
  assign _03634_ = _03633_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6303" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[10];
  assign _03635_ = _03634_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6304" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[11];
  assign _03636_ = _03635_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6304" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[12];
  assign _03637_ = _03636_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6305" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[13];
  assign _03638_ = _03637_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6305" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[14];
  assign _03639_ = _03638_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6306" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[15];
  assign _03640_ = _03639_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6306" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[16];
  assign _03641_ = _03640_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6307" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[17];
  assign _03642_ = _03641_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6307" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[18];
  assign _03643_ = _03642_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6308" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[19];
  assign _03644_ = _03643_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6308" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[20];
  assign _03645_ = _03644_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6309" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[21];
  assign _03646_ = _03645_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6309" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[22];
  assign _03647_ = _03646_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6310" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[23];
  assign _03648_ = _03647_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6310" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[25];
  assign _03649_ = FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6319" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[1];
  assign _03650_ = _03649_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6319" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[2];
  assign _03651_ = _03650_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6320" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[3];
  assign _03652_ = _03651_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6320" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[4];
  assign _03653_ = _03652_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6321" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[5];
  assign _03654_ = _03653_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6321" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[6];
  assign _03655_ = _03654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6322" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[7];
  assign _03656_ = _03655_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6322" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[8];
  assign _03657_ = _03656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6323" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[9];
  assign _03658_ = _03657_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6323" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[10];
  assign _03659_ = _03658_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6324" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[11];
  assign _03660_ = _03659_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6324" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[12];
  assign _03661_ = _03660_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6325" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[13];
  assign _03662_ = _03661_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6325" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[14];
  assign _03663_ = _03662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6326" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[15];
  assign _03664_ = _03663_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6326" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[16];
  assign _03665_ = _03664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6327" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[17];
  assign _03666_ = _03665_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6327" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[18];
  assign _03667_ = _03666_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6328" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[19];
  assign _03668_ = _03667_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6328" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[20];
  assign _03669_ = _03668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6329" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[21];
  assign _03670_ = _03669_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6329" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[22];
  assign _03671_ = _03670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6330" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[23];
  assign _03672_ = _03671_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6330" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[25];
  assign _03673_ = FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6339" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[1];
  assign _03674_ = _03673_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6339" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[2];
  assign _03675_ = _03674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6340" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[3];
  assign _03676_ = _03675_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6340" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[4];
  assign _03677_ = _03676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6341" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[5];
  assign _03678_ = _03677_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6341" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[6];
  assign _03679_ = _03678_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6342" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[7];
  assign _03680_ = _03679_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6342" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[8];
  assign _03681_ = _03680_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6343" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[9];
  assign _03682_ = _03681_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6343" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[10];
  assign _03683_ = _03682_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6344" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[11];
  assign _03684_ = _03683_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6344" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[12];
  assign _03685_ = _03684_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6345" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[13];
  assign _03686_ = _03685_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6345" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[14];
  assign _03687_ = _03686_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6346" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[15];
  assign _03688_ = _03687_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6346" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[16];
  assign _03689_ = _03688_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6347" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[17];
  assign _03690_ = _03689_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6347" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[18];
  assign _03691_ = _03690_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6348" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[19];
  assign _03692_ = _03691_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6348" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[20];
  assign _03693_ = _03692_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6349" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[21];
  assign _03694_ = _03693_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6349" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[22];
  assign _03695_ = _03694_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6350" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[23];
  assign _03696_ = _03695_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6350" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[25];
  assign _03697_ = and_1142_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6358" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp;
  assign lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1 = _03697_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6358" *) FpAdd_8U_23U_1_mux_13_itm_4;
  assign _03698_ = _02060_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6368" *) _02066_;
  assign _03699_ = IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_1_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6374" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp;
  assign lut_lookup_else_if_lor_6_lpi_1_dfm_mx0w1 = _03699_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6374" *) FpAdd_8U_23U_1_mux_29_itm_4;
  assign _03700_ = _02061_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6381" *) _02067_;
  assign _03701_ = IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_2_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6389" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp;
  assign lut_lookup_else_if_lor_7_lpi_1_dfm_mx0w1 = _03701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6389" *) FpAdd_8U_23U_1_mux_45_itm_4;
  assign _03702_ = _02062_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6396" *) _02068_;
  assign lut_lookup_if_1_lor_7_lpi_1_dfm_mx0w0 = or_2025_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6398" *) FpAdd_8U_23U_2_mux_45_itm_3;
  assign _03703_ = IsNaN_8U_23U_5_IsNaN_8U_23U_5_IsNaN_8U_23U_5_and_3_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6404" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp;
  assign lut_lookup_else_if_lor_1_lpi_1_dfm_mx0w1 = _03703_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6404" *) FpAdd_8U_23U_1_mux_61_itm_4;
  assign _03704_ = _02063_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6411" *) _02069_;
  assign lut_lookup_if_1_lor_1_lpi_1_dfm_mx0w0 = or_2035_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6413" *) FpAdd_8U_23U_2_mux_61_itm_3;
  assign lut_lookup_if_else_lut_lookup_if_else_or_3_cse = lut_lookup_if_else_else_slc_10_mdf_sva_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6416" *) _02407_;
  assign lut_lookup_if_if_lut_lookup_if_if_or_3_nl = lut_lookup_4_if_if_else_acc_nl[9] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6418" *) lut_lookup_if_if_lor_1_lpi_1_dfm_4;
  assign lut_lookup_if_else_lut_lookup_if_else_or_2_cse = lut_lookup_if_else_else_slc_10_mdf_3_sva_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6422" *) _02408_;
  assign lut_lookup_if_if_lut_lookup_if_if_or_2_nl = lut_lookup_3_if_if_else_acc_nl[9] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6424" *) lut_lookup_if_if_lor_7_lpi_1_dfm_4;
  assign lut_lookup_if_else_lut_lookup_if_else_or_1_cse = lut_lookup_if_else_else_slc_10_mdf_2_sva_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6428" *) _02409_;
  assign lut_lookup_if_if_lut_lookup_if_if_or_1_nl = lut_lookup_2_if_if_else_acc_nl[9] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6430" *) lut_lookup_if_if_lor_6_lpi_1_dfm_4;
  assign lut_lookup_if_else_lut_lookup_if_else_or_cse = lut_lookup_if_else_else_slc_10_mdf_1_sva_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6434" *) _02410_;
  assign lut_lookup_if_if_lut_lookup_if_if_or_nl = lut_lookup_1_if_if_else_acc_nl[9] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6436" *) lut_lookup_if_if_lor_5_lpi_1_dfm_4;
  assign _03705_ = _02411_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6477" *) _02071_;
  assign _03706_ = _02412_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6478" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_10_tmp;
  assign lut_lookup_if_if_lor_1_lpi_1_dfm_mx0w3 = _03706_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6478" *) FpAdd_8U_23U_1_mux_61_itm_4;
  assign _03707_ = _02413_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6483" *) _02073_;
  assign _03708_ = _02414_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6484" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_8_tmp;
  assign lut_lookup_if_if_lor_7_lpi_1_dfm_mx0w3 = _03708_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6484" *) FpAdd_8U_23U_1_mux_45_itm_4;
  assign _03709_ = _02415_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6486" *) _02075_;
  assign _03710_ = _02416_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6487" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_6_tmp;
  assign lut_lookup_if_if_lor_6_lpi_1_dfm_mx0w3 = _03710_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6487" *) FpAdd_8U_23U_1_mux_29_itm_4;
  assign _03711_ = nor_832_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6489" *) IsZero_8U_23U_5_IsZero_8U_23U_5_nor_4_tmp;
  assign lut_lookup_if_if_lor_5_lpi_1_dfm_mx0w3 = _03711_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6489" *) FpAdd_8U_23U_1_mux_13_itm_4;
  assign _03712_ = IsNaN_8U_23U_4_nor_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6549" *) IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_mx0w0;
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_4_nl = FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6587" *) _02417_;
  assign _03713_ = FpAdd_8U_23U_1_and_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6595" *) FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0;
  assign _03714_ = IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6609" *) IsNaN_8U_23U_3_land_1_lpi_1_dfm_6;
  assign FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_4_nl = FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6615" *) _02420_;
  assign _03715_ = FpAdd_8U_23U_2_and_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6623" *) FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0;
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_5_nl = FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6638" *) _02423_;
  assign _03716_ = FpAdd_8U_23U_1_and_1_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6646" *) FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0;
  assign _03717_ = IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6660" *) IsNaN_8U_23U_3_land_2_lpi_1_dfm_7;
  assign FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_5_nl = FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6668" *) _02426_;
  assign _03718_ = FpAdd_8U_23U_2_and_1_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6676" *) FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0;
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_6_nl = FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6691" *) _02429_;
  assign _03719_ = FpAdd_8U_23U_1_and_2_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6699" *) FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0;
  assign _03720_ = IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6713" *) IsNaN_8U_23U_3_land_3_lpi_1_dfm_7;
  assign FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_6_nl = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6719" *) _02432_;
  assign _03721_ = FpAdd_8U_23U_2_and_2_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6727" *) FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0;
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_7_nl = FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6742" *) _02435_;
  assign _03722_ = FpAdd_8U_23U_1_and_3_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6750" *) FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0;
  assign _03723_ = IsNaN_8U_23U_1_land_lpi_1_dfm_8 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6764" *) IsNaN_8U_23U_3_land_lpi_1_dfm_6;
  assign FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_7_nl = FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6770" *) _02438_;
  assign _03724_ = FpAdd_8U_23U_2_and_3_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6778" *) FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0;
  assign lut_lookup_lo_miss_1_sva = lut_lookup_lo_uflow_1_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6844" *) lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0;
  assign lut_lookup_le_miss_1_sva = lut_lookup_le_uflow_1_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6857" *) lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0;
  assign _03725_ = lut_lookup_le_miss_1_sva | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6867" *) lut_lookup_lo_miss_1_sva;
  assign lut_lookup_lo_miss_2_sva = lut_lookup_lo_uflow_2_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6902" *) lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0;
  assign lut_lookup_le_miss_2_sva = lut_lookup_le_uflow_2_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6903" *) lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0;
  assign _03726_ = lut_lookup_le_miss_2_sva | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6925" *) lut_lookup_lo_miss_2_sva;
  assign lut_lookup_lo_miss_3_sva = lut_lookup_lo_uflow_3_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6960" *) lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0;
  assign lut_lookup_le_miss_3_sva = lut_lookup_le_uflow_3_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6961" *) lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0;
  assign _03727_ = lut_lookup_le_miss_3_sva | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6983" *) lut_lookup_lo_miss_3_sva;
  assign lut_lookup_lo_miss_sva = lut_lookup_lo_uflow_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7018" *) lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0;
  assign lut_lookup_le_miss_sva = lut_lookup_le_uflow_lpi_1_dfm_6 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7019" *) lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0;
  assign _03728_ = lut_lookup_le_miss_sva | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7041" *) lut_lookup_lo_miss_sva;
  assign _03729_ = reg_lut_lookup_if_unequal_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7073" *) cfg_lut_le_function_1_sva_10;
  assign lut_lookup_not_39_nl = _03729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7073" *) lut_lookup_or_3_tmp;
  assign _03730_ = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7081" *) lut_lookup_1_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  assign _03731_ = _01654_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7083" *) _01655_;
  assign _03732_ = lut_lookup_1_else_2_and_svs | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7084" *) lut_lookup_1_and_svs_2;
  assign _03733_ = _01656_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7085" *) _01658_;
  assign lut_lookup_or_3_tmp = _03733_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7085" *) _01659_;
  assign lut_lookup_not_38_nl = _03729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7087" *) lut_lookup_or_7_tmp;
  assign _03734_ = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7095" *) lut_lookup_2_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  assign _03735_ = _01662_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7097" *) _01663_;
  assign _03736_ = lut_lookup_2_else_2_and_svs | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7098" *) lut_lookup_2_and_svs_2;
  assign _03737_ = _01664_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7099" *) _01666_;
  assign lut_lookup_or_7_tmp = _03737_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7099" *) _01667_;
  assign lut_lookup_not_37_nl = _03729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7101" *) lut_lookup_or_11_tmp;
  assign _03738_ = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7109" *) lut_lookup_3_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  assign _03739_ = _01668_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7111" *) _01669_;
  assign _03740_ = lut_lookup_3_else_2_and_svs | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7112" *) lut_lookup_3_and_svs_2;
  assign _03741_ = _01670_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7113" *) _01672_;
  assign lut_lookup_or_11_tmp = _03741_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7113" *) _01673_;
  assign lut_lookup_not_36_nl = _03729_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7115" *) lut_lookup_or_15_tmp;
  assign _03742_ = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7123" *) lut_lookup_4_else_2_else_lut_lookup_else_2_else_if_nor_svs;
  assign _03743_ = _01674_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7125" *) _01675_;
  assign _03744_ = lut_lookup_4_else_2_and_svs | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7126" *) lut_lookup_4_and_svs_2;
  assign _03745_ = _01676_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7127" *) _01678_;
  assign lut_lookup_or_15_tmp = _03745_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7127" *) _01679_;
  assign _03746_ = _02058_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7456" *) _02090_;
  assign _03747_ = _02074_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7458" *) _02091_;
  assign _03748_ = _02072_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7460" *) _02092_;
  assign _03749_ = _02070_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7462" *) _02093_;
  assign _03750_ = nor_874_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7464" *) _02280_;
  assign or_4_nl = _03750_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7464" *) or_1495_cse;
  assign or_tmp_8 = reg_cfg_precision_1_sva_st_12_cse_1[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7468" *) _02477_;
  assign _03751_ = or_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7472" *) _00000_;
  assign _03752_ = _03751_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7472" *) or_66_cse;
  assign or_tmp_44 = reg_cfg_precision_1_sva_st_13_cse_1[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7478" *) _02478_;
  assign _03753_ = nor_13_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7484" *) or_66_cse;
  assign or_tmp_101 = _03753_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7485" *) _00000_;
  assign _03754_ = or_66_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7490" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_6;
  assign or_tmp_124 = _03754_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7490" *) _02479_;
  assign or_122_nl = or_66_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7492" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_6;
  assign or_121_nl = or_66_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7495" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_6;
  assign _03755_ = or_1857_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7498" *) IsNaN_8U_23U_7_land_lpi_1_dfm_7;
  assign or_tmp_129 = _03755_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7498" *) _02480_;
  assign or_127_nl = or_1857_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7500" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_7;
  assign or_126_nl = or_1857_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7503" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_7;
  assign _03756_ = _03389_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7511" *) lut_lookup_2_FpMantRNE_49U_24U_2_else_and_tmp;
  assign _03757_ = _02481_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7511" *) _00000_;
  assign or_191_nl = _03757_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7511" *) or_66_cse;
  assign nand_tmp_4 = nor_874_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7514" *) mux_tmp_128;
  assign _03758_ = FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7524" *) IsNaN_8U_23U_8_land_lpi_1_dfm_5;
  assign _03759_ = _03758_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7524" *) IsNaN_8U_23U_7_land_lpi_1_dfm_7;
  assign _03760_ = _03759_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7524" *) or_1857_cse;
  assign or_302_nl = _03760_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7525" *) _00001_;
  assign _03761_ = or_969_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7532" *) _00001_;
  assign or_tmp_331 = _03761_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7532" *) or_1857_cse;
  assign _03762_ = or_1857_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7536" *) and_1140_cse;
  assign _03763_ = _03762_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7537" *) IsZero_8U_23U_8_IsZero_8U_23U_8_nor_1_tmp;
  assign _03764_ = _03763_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7537" *) FpAdd_8U_23U_2_mux_29_itm_3;
  assign or_tmp_363 = _03764_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7537" *) _00001_;
  assign or_tmp_378 = lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7540" *) not_tmp_235;
  assign _03765_ = _02978_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7543" *) or_1857_cse;
  assign or_tmp_395 = _03765_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7543" *) _00001_;
  assign _03766_ = lut_lookup_if_1_lor_7_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7544" *) _00032_;
  assign or_tmp_397 = _03766_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7544" *) or_tmp_314;
  assign _03767_ = _02975_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7548" *) or_1857_cse;
  assign or_tmp_427 = _03767_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7548" *) _00001_;
  assign _03768_ = lut_lookup_if_1_lor_1_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7549" *) _00032_;
  assign or_tmp_428 = _03768_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7549" *) or_tmp_314;
  assign _03769_ = lut_lookup_unequal_tmp_13 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7551" *) _02208_;
  assign _03770_ = _01701_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7553" *) lut_lookup_else_if_lor_5_lpi_1_dfm_st_3;
  assign _03771_ = _03770_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7553" *) _02056_;
  assign or_tmp_447 = _03771_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7553" *) _02203_;
  assign or_tmp_456 = _02056_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7555" *) _02203_;
  assign _03772_ = IsNaN_8U_23U_10_land_1_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7557" *) lut_lookup_if_1_lor_5_lpi_1_dfm_4;
  assign _03773_ = _03772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7557" *) _00032_;
  assign mux_tmp_279 = _03773_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7557" *) or_tmp_314;
  assign or_tmp_478 = _02057_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7559" *) _00010_;
  assign or_tmp_505 = cfg_precision_1_sva_st_72[0] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7564" *) not_tmp_276;
  assign _03774_ = _01704_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7566" *) lut_lookup_if_1_lor_6_lpi_1_dfm_st_4;
  assign _03775_ = _03774_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7567" *) _02057_;
  assign or_tmp_522 = _03775_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7567" *) _00010_;
  assign _03776_ = IsNaN_8U_23U_10_land_2_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7569" *) lut_lookup_if_1_lor_6_lpi_1_dfm_4;
  assign _03777_ = _03776_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7569" *) _00032_;
  assign mux_tmp_301 = _03777_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7569" *) or_tmp_314;
  assign _03778_ = _01705_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7572" *) lut_lookup_else_if_lor_7_lpi_1_dfm_st_3;
  assign _03779_ = _03778_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7572" *) _02056_;
  assign or_tmp_547 = _03779_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7572" *) _02203_;
  assign _03780_ = IsNaN_8U_23U_10_land_3_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7575" *) lut_lookup_if_1_lor_7_lpi_1_dfm_4;
  assign _03781_ = _03780_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7575" *) _00032_;
  assign or_tmp_573 = _03781_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7575" *) or_tmp_314;
  assign _03782_ = _01706_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7577" *) lut_lookup_else_if_lor_1_lpi_1_dfm_st_3;
  assign _03783_ = _03782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7577" *) _02056_;
  assign or_tmp_598 = _03783_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7577" *) _02203_;
  assign _03784_ = IsNaN_8U_23U_10_land_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7580" *) lut_lookup_if_1_lor_1_lpi_1_dfm_4;
  assign _03785_ = _03784_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7580" *) _00032_;
  assign or_tmp_623 = _03785_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7580" *) or_tmp_314;
  assign _03786_ = cfg_lut_le_function_1_sva_10 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7581" *) _00010_;
  assign _03787_ = reg_cfg_precision_1_sva_st_12_cse_1[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7584" *) _02482_;
  assign _00016_ = reg_cfg_precision_1_sva_st_12_cse_1[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7585" *) or_1689_cse;
  assign _03788_ = reg_cfg_precision_1_sva_st_12_cse_1[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7586" *) _00003_;
  assign _03789_ = reg_cfg_precision_1_sva_st_12_cse_1[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7587" *) _00033_;
  assign _03790_ = IsNaN_8U_23U_8_land_2_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7595" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
  assign _03791_ = _03790_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7595" *) _00033_;
  assign or_1860_nl = _03791_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7595" *) mux_tmp_595;
  assign or_tmp_843 = or_1495_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7597" *) _02483_;
  assign or_841_nl = _00000_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7601" *) reg_cfg_precision_1_sva_st_13_cse_1[0];
  assign _03792_ = lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7604" *) _02484_;
  assign or_832_nl = IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7605" *) IsNaN_8U_23U_8_land_2_lpi_1_dfm_5;
  assign _03793_ = reg_cfg_precision_1_sva_st_13_cse_1[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7613" *) _00000_;
  assign _03794_ = cfg_precision_1_sva_st_70[1] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7616" *) _00001_;
  assign _03795_ = or_1857_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7620" *) cfg_lut_le_function_1_sva_st_41;
  assign or_tmp_976 = _03795_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7620" *) _00001_;
  assign _03796_ = or_1202_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7622" *) cfg_lut_le_function_1_sva_st_42;
  assign or_tmp_980 = _03796_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7622" *) _00032_;
  assign _03797_ = nor_610_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7623" *) cfg_lut_le_function_1_sva_st_42;
  assign or_tmp_993 = _03797_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7623" *) _00032_;
  assign _03798_ = FpMantRNE_49U_24U_2_else_carry_1_sva_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7633" *) FpAdd_8U_23U_2_mux_13_itm_3;
  assign or_tmp_1043 = _03798_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7633" *) _02485_;
  assign _03799_ = nor_792_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *) FpMantRNE_49U_24U_2_else_carry_2_sva_2;
  assign _03800_ = _03799_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *) FpAdd_8U_23U_2_mux_29_itm_3;
  assign _03801_ = _03800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7642" *) _02486_;
  assign _03802_ = FpAdd_8U_23U_2_mux_45_itm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7651" *) _02269_;
  assign _03803_ = _03802_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7651" *) FpMantRNE_49U_24U_2_else_carry_3_sva_2;
  assign or_tmp_1181 = _03803_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7652" *) _02488_;
  assign _03804_ = FpMantRNE_49U_24U_2_else_carry_sva_2 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7661" *) FpAdd_8U_23U_2_mux_61_itm_3;
  assign or_tmp_1250 = _03804_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7661" *) _02489_;
  assign _03805_ = and_794_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7665" *) _02280_;
  assign or_tmp_1360 = _03805_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7665" *) or_1495_cse;
  assign _03806_ = or_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7669" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign or_tmp_1450 = _03806_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7669" *) not_tmp_800;
  assign or_tmp_1490 = or_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7682" *) or_66_cse;
  assign or_dcpl_51 = nor_193_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7685" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign or_dcpl_57 = and_dcpl_98 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7688" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _03807_ = _02491_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7690" *) IsNaN_8U_23U_6_land_1_lpi_1_dfm_6;
  assign _03808_ = _03807_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7690" *) or_tmp_314;
  assign or_1583_nl = lut_lookup_if_if_lor_5_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7690" *) _02492_;
  assign or_tmp_1513 = lut_lookup_lo_uflow_1_lpi_1_dfm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7694" *) mux_tmp_1130;
  assign _03809_ = _02493_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7697" *) IsNaN_8U_23U_6_land_2_lpi_1_dfm_6;
  assign _03810_ = _03809_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7697" *) or_tmp_314;
  assign or_1594_nl = lut_lookup_if_if_lor_6_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7697" *) _02494_;
  assign or_tmp_1523 = lut_lookup_lo_uflow_2_lpi_1_dfm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7702" *) mux_tmp_1143;
  assign _03811_ = _02495_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7705" *) IsNaN_8U_23U_6_land_3_lpi_1_dfm_6;
  assign _03812_ = _03811_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7705" *) or_tmp_314;
  assign or_1606_nl = lut_lookup_if_if_lor_7_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7705" *) _02496_;
  assign or_tmp_1534 = lut_lookup_lo_uflow_3_lpi_1_dfm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7710" *) mux_tmp_1156;
  assign _03813_ = _02497_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7713" *) IsNaN_8U_23U_6_land_lpi_1_dfm_6;
  assign _03814_ = _03813_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7713" *) or_tmp_314;
  assign or_1618_nl = lut_lookup_if_if_lor_1_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7713" *) _02498_;
  assign or_tmp_1545 = lut_lookup_lo_uflow_lpi_1_dfm_3 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7718" *) mux_tmp_1169;
  assign _03815_ = _02500_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7723" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl[23];
  assign _03816_ = _02501_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7725" *) FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl[23];
  assign _03817_ = _02503_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7727" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl[23];
  assign _03818_ = _02505_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7729" *) FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl[23];
  assign _03819_ = _02507_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7731" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl[23];
  assign _03820_ = _02509_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7733" *) FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl[23];
  assign _03821_ = _02512_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7735" *) FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl[23];
  assign _03822_ = _02513_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7737" *) FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl[23];
  assign chn_lut_in_rsci_ld_core_psct_mx0c0 = main_stage_en_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7747" *) fsm_output[0];
  assign _03823_ = cfg_lut_uflow_priority_1_sva_9 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7754" *) _02516_;
  assign _03824_ = cfg_lut_uflow_priority_1_sva_9 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7759" *) _02517_;
  assign _03825_ = cfg_lut_uflow_priority_1_sva_9 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7764" *) _02518_;
  assign _03826_ = cfg_lut_uflow_priority_1_sva_9 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7769" *) _02519_;
  assign _03827_ = IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7814" *) reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign _03828_ = reg_cfg_lut_le_function_1_sva_st_19_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7817" *) reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse;
  assign _03829_ = nor_193_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7822" *) _00000_;
  assign _03830_ = _03829_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7823" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _03831_ = _03830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7823" *) lut_lookup_1_if_else_else_acc_nl[10];
  assign or_tmp_1663 = _03831_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7823" *) _02530_;
  assign or_tmp_1671 = _02530_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7825" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _03832_ = _03830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7827" *) lut_lookup_2_if_else_else_acc_nl[10];
  assign or_tmp_1674 = _03832_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7827" *) _02173_;
  assign or_tmp_1678 = or_40_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7829" *) lut_lookup_2_if_else_else_acc_nl[10];
  assign _03833_ = _03830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7831" *) lut_lookup_3_if_else_else_acc_nl[10];
  assign or_tmp_1684 = _03833_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7831" *) _02343_;
  assign or_1972_nl = IsNaN_8U_23U_4_land_3_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7832" *) nor_38_cse_1;
  assign or_1973_nl = IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7833" *) nor_38_cse_1;
  assign _03834_ = IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7836" *) mux_1234_nl;
  assign or_tmp_1692 = lut_lookup_3_FpMantRNE_49U_24U_else_and_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7836" *) _02531_;
  assign _03835_ = _03830_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7838" *) lut_lookup_4_if_else_else_acc_nl[10];
  assign or_tmp_1697 = _03835_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7838" *) _02532_;
  assign or_1991_nl = IsNaN_8U_23U_4_land_lpi_1_dfm_4 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7839" *) nor_50_cse_1;
  assign or_1992_nl = reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7840" *) nor_50_cse_1;
  assign _03836_ = IsNaN_8U_23U_1_land_lpi_1_dfm_7 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7843" *) mux_1241_nl;
  assign or_tmp_1705 = lut_lookup_4_FpMantRNE_49U_24U_else_and_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7843" *) _02533_;
  assign or_tmp_1707 = _02532_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7844" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _03837_ = _02258_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7847" *) FpMantRNE_49U_24U_2_else_carry_1_sva_2;
  assign or_tmp_1716 = _03837_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7847" *) _02096_;
  assign _03838_ = nor_792_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7848" *) _02264_;
  assign _03839_ = _03838_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7849" *) FpMantRNE_49U_24U_2_else_carry_2_sva_2;
  assign or_tmp_1720 = _03839_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7849" *) _02097_;
  assign _03840_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7851" *) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247];
  assign _03841_ = _02534_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7852" *) lut_lookup_if_1_lor_5_lpi_1_dfm_5;
  assign _03842_ = _03841_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7852" *) IsNaN_8U_23U_10_land_1_lpi_1_dfm_6;
  assign _03843_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7856" *) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247];
  assign _03844_ = lut_lookup_if_1_lor_6_lpi_1_dfm_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7856" *) _02535_;
  assign _03845_ = _03844_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7856" *) IsNaN_8U_23U_10_land_2_lpi_1_dfm_6;
  assign _03846_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7860" *) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247];
  assign _03847_ = _02536_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7861" *) lut_lookup_if_1_lor_7_lpi_1_dfm_5;
  assign _03848_ = _03847_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7861" *) IsNaN_8U_23U_10_land_3_lpi_1_dfm_6;
  assign _03849_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7864" *) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247];
  assign or_2056_nl = lut_lookup_unequal_tmp_13 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7865" *) _00087_[34];
  assign or_2055_nl = nor_813_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7866" *) lut_lookup_if_1_lor_1_lpi_1_dfm_5;
  assign _03850_ = or_2055_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7869" *) lut_lookup_unequal_tmp_13;
  assign _03851_ = _03850_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7869" *) IsNaN_8U_23U_10_land_lpi_1_dfm_6;
  assign _03852_ = and_dcpl_72 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8086" *) and_dcpl_74;
  assign _03853_ = or_tmp_1628 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8094" *) main_stage_v_1_mx0c1;
  assign _03854_ = IsNaN_8U_23U_3_nor_10_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8197" *) _02094_;
  assign _03855_ = IsNaN_8U_23U_3_nor_4_tmp | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8211" *) _02095_;
  assign _03856_ = IsNaN_8U_23U_8_nor_2_tmp_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8217" *) IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_mx0w0;
  assign _03857_ = _01782_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8224" *) main_stage_v_2_mx0c1;
  assign _03858_ = and_956_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8278" *) _01787_;
  assign _03859_ = and_284_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8286" *) and_286_rgt;
  assign _03860_ = _03859_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8286" *) and_288_rgt;
  assign _03861_ = _03860_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8286" *) and_290_rgt;
  assign _03862_ = _01792_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8311" *) and_292_rgt;
  assign _03863_ = and_956_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8333" *) _01795_;
  assign _03864_ = and_300_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8341" *) and_302_rgt;
  assign _03865_ = _03864_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8341" *) and_304_rgt;
  assign _03866_ = _03865_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8341" *) and_306_rgt;
  assign _03867_ = _01800_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8364" *) and_308_rgt;
  assign _03868_ = and_956_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8373" *) _01803_;
  assign _03869_ = and_316_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8382" *) and_318_rgt;
  assign _03870_ = _03869_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8382" *) and_320_rgt;
  assign _03871_ = _03870_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8382" *) and_322_rgt;
  assign _03872_ = _01808_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8413" *) and_324_rgt;
  assign _03873_ = and_956_cse | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8422" *) _01811_;
  assign _03874_ = and_330_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8431" *) and_332_rgt;
  assign _03875_ = _03874_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8431" *) and_334_rgt;
  assign _03876_ = _03875_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8431" *) and_336_rgt;
  assign _03877_ = _01816_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8444" *) and_338_rgt;
  assign _03878_ = _01819_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8453" *) main_stage_v_3_mx0c1;
  assign _03879_ = and_344_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8503" *) and_dcpl_148;
  assign _03880_ = _03879_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8503" *) and_347_rgt;
  assign _03881_ = lut_lookup_1_if_else_else_acc_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8526" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _03882_ = FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8676" *) FpAdd_8U_23U_2_and_4_rgt;
  assign _03883_ = _03882_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8676" *) FpAdd_8U_23U_2_and_5_rgt;
  assign _03884_ = lut_lookup_2_if_else_else_acc_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8746" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _03885_ = FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_1_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8835" *) FpAdd_8U_23U_2_and_10_rgt;
  assign _03886_ = _03885_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8835" *) FpAdd_8U_23U_2_and_11_rgt;
  assign _03887_ = lut_lookup_3_if_else_else_acc_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8894" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _03888_ = mux_1233_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8915" *) nor_38_cse_1;
  assign _03889_ = _03888_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8915" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign _03890_ = _02571_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8916" *) lut_lookup_3_FpMantRNE_49U_24U_else_and_tmp;
  assign _03891_ = FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_2_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8969" *) FpAdd_8U_23U_2_and_16_rgt;
  assign _03892_ = _03891_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8969" *) FpAdd_8U_23U_2_and_17_rgt;
  assign _03893_ = lut_lookup_4_if_else_else_acc_nl[10] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9014" *) reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _03894_ = mux_1240_nl | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9035" *) nor_50_cse_1;
  assign _03895_ = _03894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9035" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _03896_ = _02577_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9036" *) lut_lookup_4_FpMantRNE_49U_24U_else_and_tmp;
  assign _03897_ = FpAdd_8U_23U_2_o_expo_FpAdd_8U_23U_2_o_expo_nor_3_rgt | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9089" *) FpAdd_8U_23U_2_and_22_rgt;
  assign _03898_ = _03897_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9089" *) FpAdd_8U_23U_2_and_23_rgt;
  assign _03899_ = _01894_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9111" *) main_stage_v_4_mx0c1;
  assign _03900_ = _01925_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9433" *) main_stage_v_5_mx0c1;
  assign _03901_ = _01983_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9589" *) lut_lookup_else_2_else_else_if_mux_5_itm_1_mx0c1;
  assign _03902_ = _01995_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9719" *) lut_lookup_else_2_else_else_if_mux_12_itm_1_mx0c1;
  assign _03903_ = _02007_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9813" *) lut_lookup_else_2_else_else_if_mux_19_itm_1_mx0c1;
  assign _03904_ = _02017_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9911" *) lut_lookup_else_2_else_else_if_mux_26_itm_1_mx0c1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_1_sva_5 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_1_sva_5 <= _00471_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_sva_5 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_sva_5 <= _00483_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_3_sva_5 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_3_sva_5 <= _00479_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_2_sva_5 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_2_sva_5 <= _00475_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_sva_6 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_sva_6 <= _00484_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_le_data_sub_sva_1_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      lut_lookup_if_else_else_le_data_sub_sva_1_30_0_1 <= _00569_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_le_data_sub_3_sva_1_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      lut_lookup_if_else_else_le_data_sub_3_sva_1_30_0_1 <= _00568_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_3_sva_6 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_3_sva_6 <= _00480_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_2_sva_6 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_2_sva_6 <= _00476_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_le_data_sub_2_sva_1_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      lut_lookup_if_else_else_le_data_sub_2_sva_1_30_0_1 <= _00567_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_1_sva_6 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_1_sva_6 <= _00472_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_le_data_sub_1_sva_1_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      lut_lookup_if_else_else_le_data_sub_1_sva_1_30_0_1 <= _00566_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lo_index_u_sva_4 <= 32'd0;
    else
      lut_lookup_else_1_lo_index_u_sva_4 <= _00466_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_le_index_u_sva_4 <= 32'd0;
    else
      lut_lookup_else_else_else_le_index_u_sva_4 <= _00510_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 <= 6'b000000;
    else
      lut_lookup_4_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 <= _00453_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lo_index_u_3_sva_4 <= 32'd0;
    else
      lut_lookup_else_1_lo_index_u_3_sva_4 <= _00464_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_le_index_u_3_sva_4 <= 32'd0;
    else
      lut_lookup_else_else_else_le_index_u_3_sva_4 <= _00508_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 <= 6'b000000;
    else
      lut_lookup_3_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 <= _00427_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lo_index_u_2_sva_4 <= 32'd0;
    else
      lut_lookup_else_1_lo_index_u_2_sva_4 <= _00462_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_le_index_u_2_sva_4 <= 32'd0;
    else
      lut_lookup_else_else_else_le_index_u_2_sva_4 <= _00506_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 <= 6'b000000;
    else
      lut_lookup_2_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 <= _00402_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lo_index_u_1_sva_4 <= 32'd0;
    else
      lut_lookup_else_1_lo_index_u_1_sva_4 <= _00460_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_le_index_u_1_sva_4 <= 32'd0;
    else
      lut_lookup_else_else_else_le_index_u_1_sva_4 <= _00504_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 <= 6'b000000;
    else
      lut_lookup_1_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 <= _00377_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_8_nor_3_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_8_nor_3_itm_2 <= _00265_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_3_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_3_itm_2 <= _00256_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_49_itm_2 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_49_itm_2 <= _00147_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2 <= _00222_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_4_nor_3_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_4_nor_3_itm_2 <= _00228_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_49_itm_2 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_49_itm_2 <= _00115_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_8_nor_2_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_8_nor_2_itm_2 <= _00264_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_2 <= _00255_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_33_itm_2 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_33_itm_2 <= _00144_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_33_itm_2 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_33_itm_2 <= _00112_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_17_itm_2 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_17_itm_2 <= _00140_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_17_itm_2 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_17_itm_2 <= _00108_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_1_itm_2 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_1_itm_2 <= _00141_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2 <= _00223_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_4_nor_itm_2 <= 1'b0;
    else
      IsNaN_8U_23U_4_nor_itm_2 <= _00229_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_1_itm_2 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_1_itm_2 <= _00109_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_11 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_11 <= _00635_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_11 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_11 <= _00632_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_11 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_11 <= _00629_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_11 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_11 <= _00626_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 <= 1'b0;
    else
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 <= _00371_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 <= 1'b0;
    else
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 <= _00396_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 <= 1'b0;
    else
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 <= _00421_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 <= 1'b0;
    else
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 <= _00447_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_1_sva_7 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_1_sva_7 <= _00473_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_3_sva_7 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_3_sva_7 <= _00481_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_2_sva_7 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_2_sva_7 <= _00477_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_sva_7 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_sva_7 <= _00485_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_sva_3 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_sva_3 <= _00500_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntLog2_32U_ac_int_cctor_1_30_0_sva_1 <= 31'b0000000000000000000000000000000;
    else
      IntLog2_32U_ac_int_cctor_1_30_0_sva_1 <= _00193_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_3_sva_3 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_3_sva_3 <= _00497_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntLog2_32U_ac_int_cctor_1_30_0_3_sva_1 <= 31'b0000000000000000000000000000000;
    else
      IntLog2_32U_ac_int_cctor_1_30_0_3_sva_1 <= _00192_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_2_sva_3 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_2_sva_3 <= _00494_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_slc_32_mdf_sva_7 <= 1'b0;
    else
      lut_lookup_else_else_slc_32_mdf_sva_7 <= _00521_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_slc_32_mdf_3_sva_7 <= 1'b0;
    else
      lut_lookup_else_else_slc_32_mdf_3_sva_7 <= _00519_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_slc_32_mdf_2_sva_7 <= 1'b0;
    else
      lut_lookup_else_else_slc_32_mdf_2_sva_7 <= _00517_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntLog2_32U_ac_int_cctor_1_30_0_2_sva_1 <= 31'b0000000000000000000000000000000;
    else
      IntLog2_32U_ac_int_cctor_1_30_0_2_sva_1 <= _00191_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_1_sva_3 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_1_sva_3 <= _00491_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_slc_32_mdf_1_sva_7 <= 1'b0;
    else
      lut_lookup_else_else_slc_32_mdf_1_sva_7 <= _00515_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IntLog2_32U_ac_int_cctor_1_30_0_1_sva_2 <= 31'b0000000000000000000000000000000;
    else
      IntLog2_32U_ac_int_cctor_1_30_0_1_sva_2 <= _00190_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_mux_itm_2 <= 1'b0;
    else
      lut_lookup_else_mux_itm_2 <= _00542_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_mux_43_itm_2 <= 1'b0;
    else
      lut_lookup_else_mux_43_itm_2 <= _00540_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_mux_86_itm_2 <= 1'b0;
    else
      lut_lookup_else_mux_86_itm_2 <= _00541_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_mux_129_itm_2 <= 1'b0;
    else
      lut_lookup_else_mux_129_itm_2 <= _00539_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3 <= 1'b0;
    else
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3 <= _00450_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_4_else_1_else_else_acc_1_itm <= 8'b00000000;
    else
      reg_lut_lookup_4_else_1_else_else_acc_1_itm <= _00719_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_4_else_1_else_else_acc_itm <= 1'b0;
    else
      reg_lut_lookup_4_else_1_else_else_acc_itm <= _00720_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_else_1_else_else_lo_data_f_and_itm_2 <= 32'd0;
    else
      lut_lookup_4_else_1_else_else_lo_data_f_and_itm_2 <= _00446_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5 <= 23'b00000000000000000000000;
    else
      FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5 <= _00157_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_sva_4 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_sva_4 <= _00501_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_4_else_else_else_else_acc_2_reg <= 3'b000;
    else
      reg_lut_lookup_4_else_else_else_else_acc_2_reg <= _00722_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_else_else_else_else_le_data_f_and_itm_2 <= 32'd0;
    else
      lut_lookup_4_else_else_else_else_le_data_f_and_itm_2 <= _00451_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 <= 2'b00;
    else
      lut_lookup_4_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 <= _00444_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_if_else_slc_32_svs_8 <= 1'b0;
    else
      lut_lookup_4_if_else_slc_32_svs_8 <= _00457_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_sva_4 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_sva_4 <= _00580_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_else_asn_mdf_sva_2 <= 1'b0;
    else
      lut_lookup_if_else_else_else_asn_mdf_sva_2 <= _00565_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_if_lor_1_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_if_if_lor_1_lpi_1_dfm_4 <= _00582_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_sva_8 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_sva_8 <= _00486_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_3_sva_8 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_3_sva_8 <= _00482_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3 <= 1'b0;
    else
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3 <= _00424_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_3_else_1_else_else_acc_1_itm <= 8'b00000000;
    else
      reg_lut_lookup_3_else_1_else_else_acc_1_itm <= _00708_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_3_else_1_else_else_acc_itm <= 1'b0;
    else
      reg_lut_lookup_3_else_1_else_else_acc_itm <= _00709_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_else_1_else_else_lo_data_f_and_itm_2 <= 32'd0;
    else
      lut_lookup_3_else_1_else_else_lo_data_f_and_itm_2 <= _00420_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5 <= 23'b00000000000000000000000;
    else
      FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5 <= _00156_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_3_sva_4 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_3_sva_4 <= _00498_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_3_else_else_else_else_acc_2_reg <= 3'b000;
    else
      reg_lut_lookup_3_else_else_else_else_acc_2_reg <= _00711_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_else_else_else_else_le_data_f_and_itm_2 <= 32'd0;
    else
      lut_lookup_3_else_else_else_else_le_data_f_and_itm_2 <= _00425_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 <= 2'b00;
    else
      lut_lookup_3_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 <= _00418_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_3_sva_4 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_3_sva_4 <= _00577_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_else_asn_mdf_3_sva_2 <= 1'b0;
    else
      lut_lookup_if_else_else_else_asn_mdf_3_sva_2 <= _00564_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_2_sva_8 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_2_sva_8 <= _00478_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3 <= 1'b0;
    else
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3 <= _00399_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_2_else_1_else_else_acc_1_itm <= 8'b00000000;
    else
      reg_lut_lookup_2_else_1_else_else_acc_1_itm <= _00697_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_2_else_1_else_else_acc_itm <= 1'b0;
    else
      reg_lut_lookup_2_else_1_else_else_acc_itm <= _00698_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_else_1_else_else_lo_data_f_and_itm_2 <= 32'd0;
    else
      lut_lookup_2_else_1_else_else_lo_data_f_and_itm_2 <= _00395_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5 <= 23'b00000000000000000000000;
    else
      FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5 <= _00155_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_slc_32_mdf_sva_8 <= 1'b0;
    else
      lut_lookup_else_else_slc_32_mdf_sva_8 <= _00522_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_slc_32_mdf_3_sva_8 <= 1'b0;
    else
      lut_lookup_else_else_slc_32_mdf_3_sva_8 <= _00520_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_slc_32_mdf_2_sva_8 <= 1'b0;
    else
      lut_lookup_else_else_slc_32_mdf_2_sva_8 <= _00518_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_2_sva_4 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_2_sva_4 <= _00495_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_2_else_else_else_else_acc_2_reg <= 3'b000;
    else
      reg_lut_lookup_2_else_else_else_else_acc_2_reg <= _00700_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_else_else_else_else_le_data_f_and_itm_2 <= 32'd0;
    else
      lut_lookup_2_else_else_else_else_le_data_f_and_itm_2 <= _00400_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 <= 2'b00;
    else
      lut_lookup_2_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 <= _00393_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg <= 8'b00000000;
    else
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg <= _00671_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg <= 8'b00000000;
    else
      reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg <= _00674_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IntLog2_32U_ac_int_cctor_1_30_0_reg <= 8'b00000000;
    else
      reg_IntLog2_32U_ac_int_cctor_1_30_0_reg <= _00675_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_2_sva_4 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_2_sva_4 <= _00574_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_else_asn_mdf_2_sva_2 <= 1'b0;
    else
      lut_lookup_if_else_else_else_asn_mdf_2_sva_2 <= _00563_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_slc_32_mdf_1_sva_8 <= 1'b0;
    else
      lut_lookup_else_1_slc_32_mdf_1_sva_8 <= _00474_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3 <= 1'b0;
    else
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3 <= _00374_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_1_else_1_else_else_acc_1_itm <= 8'b00000000;
    else
      reg_lut_lookup_1_else_1_else_else_acc_1_itm <= _00686_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_1_else_1_else_else_acc_itm <= 1'b0;
    else
      reg_lut_lookup_1_else_1_else_else_acc_itm <= _00687_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_else_1_else_else_lo_data_f_and_itm_2 <= 32'd0;
    else
      lut_lookup_1_else_1_else_else_lo_data_f_and_itm_2 <= _00370_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5 <= 23'b00000000000000000000000;
    else
      FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5 <= _00154_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_slc_32_mdf_1_sva_8 <= 1'b0;
    else
      lut_lookup_else_else_slc_32_mdf_1_sva_8 <= _00516_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_1_sva_4 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_1_sva_4 <= _00492_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_1_else_else_else_else_acc_3_reg <= 4'b0000;
    else
      reg_lut_lookup_1_else_else_else_else_acc_3_reg <= _00690_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg <= 23'b00000000000000000000000;
    else
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg <= _00670_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_2_else_else_else_else_acc_3_reg <= 4'b0000;
    else
      reg_lut_lookup_2_else_else_else_else_acc_3_reg <= _00701_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg <= 23'b00000000000000000000000;
    else
      reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg <= _00673_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_3_else_else_else_else_acc_3_reg <= 4'b0000;
    else
      reg_lut_lookup_3_else_else_else_else_acc_3_reg <= _00712_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 <= 23'b00000000000000000000000;
    else
      reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 <= _00672_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_4_else_else_else_else_acc_3_reg <= 4'b0000;
    else
      reg_lut_lookup_4_else_else_else_else_acc_3_reg <= _00723_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_1_else_else_else_else_acc_2_reg <= 3'b000;
    else
      reg_lut_lookup_1_else_else_else_else_acc_2_reg <= _00689_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_1_else_else_else_else_acc_1_reg <= 1'b0;
    else
      reg_lut_lookup_1_else_else_else_else_acc_1_reg <= _00688_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_2_else_else_else_else_acc_1_reg <= 1'b0;
    else
      reg_lut_lookup_2_else_else_else_else_acc_1_reg <= _00699_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_3_else_else_else_else_acc_1_reg <= 1'b0;
    else
      reg_lut_lookup_3_else_else_else_else_acc_1_reg <= _00710_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_4_else_else_else_else_acc_1_reg <= 1'b0;
    else
      reg_lut_lookup_4_else_else_else_else_acc_1_reg <= _00721_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_1_else_else_else_else_acc_reg <= 1'b0;
    else
      reg_lut_lookup_1_else_else_else_else_acc_reg <= _00691_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_2_else_else_else_else_acc_reg <= 1'b0;
    else
      reg_lut_lookup_2_else_else_else_else_acc_reg <= _00702_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_3_else_else_else_else_acc_reg <= 1'b0;
    else
      reg_lut_lookup_3_else_else_else_else_acc_reg <= _00713_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_4_else_else_else_else_acc_reg <= 1'b0;
    else
      reg_lut_lookup_4_else_else_else_else_acc_reg <= _00724_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_else_else_else_else_le_data_f_and_itm_2 <= 32'd0;
    else
      lut_lookup_1_else_else_else_else_le_data_f_and_itm_2 <= _00375_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_precision_1_sva_8 <= 2'b00;
    else
      cfg_precision_1_sva_8 <= _00300_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 <= 2'b00;
    else
      lut_lookup_1_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 <= _00368_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm <= 23'b00000000000000000000000;
    else
      reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm <= _00668_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm <= 8'b00000000;
    else
      reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm <= _00669_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_if_else_slc_32_svs_8 <= 1'b0;
    else
      lut_lookup_3_if_else_slc_32_svs_8 <= _00431_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_if_else_slc_32_svs_8 <= 1'b0;
    else
      lut_lookup_2_if_else_slc_32_svs_8 <= _00406_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_if_else_slc_32_svs_8 <= 1'b0;
    else
      lut_lookup_1_if_else_slc_32_svs_8 <= _00381_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_1_sva_4 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_1_sva_4 <= _00571_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_else_asn_mdf_1_sva_2 <= 1'b0;
    else
      lut_lookup_if_else_else_else_asn_mdf_1_sva_2 <= _00562_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_if_lor_7_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_if_if_lor_7_lpi_1_dfm_4 <= _00585_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_if_lor_6_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_if_if_lor_6_lpi_1_dfm_4 <= _00584_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_if_lor_5_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_if_if_lor_5_lpi_1_dfm_4 <= _00583_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_10_land_1_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_8U_23U_10_land_1_lpi_1_dfm_5 <= _00194_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_6_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_if_1_lor_6_lpi_1_dfm_4 <= _00556_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_5_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_if_1_lor_5_lpi_1_dfm_4 <= _00553_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_10_land_2_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_8U_23U_10_land_2_lpi_1_dfm_5 <= _00196_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_12 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_12 <= _00630_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_12 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_12 <= _00627_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 <= 1'b0;
    else
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 <= _00372_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 <= 1'b0;
    else
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 <= _00397_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_10_land_3_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_8U_23U_10_land_3_lpi_1_dfm_5 <= _00198_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_1_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_if_1_lor_1_lpi_1_dfm_4 <= _00550_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_7_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_if_1_lor_7_lpi_1_dfm_4 <= _00559_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_10_land_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_8U_23U_10_land_lpi_1_dfm_5 <= _00200_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_12 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_12 <= _00636_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_12 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_12 <= _00633_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 <= 1'b0;
    else
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 <= _00422_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 <= 1'b0;
    else
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4 <= _00448_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_5_lpi_1_dfm_5 <= 1'b0;
    else
      lut_lookup_else_if_lor_5_lpi_1_dfm_5 <= _00530_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_6_land_1_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_6_land_1_lpi_1_dfm_6 <= _00230_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 <= _00232_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 <= _00234_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_unequal_tmp_12 <= 1'b0;
    else
      lut_lookup_else_unequal_tmp_12 <= _00543_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_1_lpi_1_dfm_5 <= 1'b0;
    else
      lut_lookup_else_if_lor_1_lpi_1_dfm_5 <= _00527_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_7_lpi_1_dfm_5 <= 1'b0;
    else
      lut_lookup_else_if_lor_7_lpi_1_dfm_5 <= _00536_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_6_lpi_1_dfm_5 <= 1'b0;
    else
      lut_lookup_else_if_lor_6_lpi_1_dfm_5 <= _00533_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_6_land_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_6_land_lpi_1_dfm_6 <= _00236_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lo_index_u_sva_3 <= 32'd0;
    else
      lut_lookup_else_1_lo_index_u_sva_3 <= _00465_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_le_index_u_sva_3 <= 32'd0;
    else
      lut_lookup_else_else_else_le_index_u_sva_3 <= _00509_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lo_index_u_3_sva_3 <= 32'd0;
    else
      lut_lookup_else_1_lo_index_u_3_sva_3 <= _00463_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_le_index_u_3_sva_3 <= 32'd0;
    else
      lut_lookup_else_else_else_le_index_u_3_sva_3 <= _00507_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lo_index_u_2_sva_3 <= 32'd0;
    else
      lut_lookup_else_1_lo_index_u_2_sva_3 <= _00461_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_le_index_u_2_sva_3 <= 32'd0;
    else
      lut_lookup_else_else_else_le_index_u_2_sva_3 <= _00505_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lo_index_u_1_sva_3 <= 32'd0;
    else
      lut_lookup_else_1_lo_index_u_1_sva_3 <= _00459_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_le_index_u_1_sva_3 <= 32'd0;
    else
      lut_lookup_else_else_else_le_index_u_1_sva_3 <= _00503_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_61_itm_1 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_61_itm_1 <= _00148_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_61_itm_3 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_61_itm_3 <= _00116_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_45_itm_1 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_45_itm_1 <= _00145_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_45_itm_3 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_45_itm_3 <= _00113_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_29_itm_1 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_29_itm_1 <= _00142_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_29_itm_3 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_29_itm_3 <= _00110_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_13_itm_1 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_13_itm_1 <= _00138_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_13_itm_3 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_13_itm_3 <= _00106_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 <= _00243_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 <= _00247_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_lpi_1_dfm_6 <= _00252_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_4_land_1_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_8U_23U_4_land_1_lpi_1_dfm_4 <= _00224_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 <= _00208_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 <= _00206_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_lpi_1_dfm_7 <= _00211_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 <= _00203_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 <= _00238_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_4_land_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_8U_23U_4_land_lpi_1_dfm_4 <= _00227_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_4_land_3_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_8U_23U_4_land_3_lpi_1_dfm_5 <= _00226_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_4_land_2_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_8U_23U_4_land_2_lpi_1_dfm_5 <= _00225_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_a_right_shift_qr_sva_3 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_a_right_shift_qr_sva_3 <= _00125_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= 1'b0;
    else
      lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= _00435_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2 <= 1'b0;
    else
      lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2 <= _00436_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_a_right_shift_qr_3_sva_3 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_a_right_shift_qr_3_sva_3 <= _00124_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= 1'b0;
    else
      lut_lookup_3_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= _00410_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_lpi_1_dfm_6 <= _00210_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
    else
      lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= _00383_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= 1'b0;
    else
      lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= _00384_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
    else
      lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= _00408_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= 1'b0;
    else
      lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= _00409_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
    else
      lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= _00433_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= 1'b0;
    else
      lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= _00434_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4 <= 1'b0;
    else
      FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4 <= _00130_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4 <= 1'b0;
    else
      FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4 <= _00131_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4 <= 1'b0;
    else
      FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4 <= _00132_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4 <= 1'b0;
    else
      FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4 <= _00133_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 <= _00202_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
    else
      lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= _00358_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= 1'b0;
    else
      lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2 <= _00359_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 <= 1'b0;
    else
      FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 <= _00098_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 <= 1'b0;
    else
      FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 <= _00099_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 <= 1'b0;
    else
      FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 <= _00100_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 <= 1'b0;
    else
      FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 <= _00101_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_qr_lpi_1_dfm_4 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_qr_lpi_1_dfm_4 <= _00164_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_qr_4_lpi_1_dfm_4 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_qr_4_lpi_1_dfm_4 <= _00162_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_a_right_shift_qr_2_sva_3 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_a_right_shift_qr_2_sva_3 <= _00123_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_qr_3_lpi_1_dfm_4 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_qr_3_lpi_1_dfm_4 <= _00160_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_a_right_shift_qr_1_sva_3 <= 8'b00000000;
    else
      FpAdd_8U_23U_1_a_right_shift_qr_1_sva_3 <= _00090_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_qr_2_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_1_qr_2_lpi_1_dfm_5 <= _00118_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_uflow_1_lpi_1_dfm_3 <= 1'b0;
    else
      lut_lookup_lo_uflow_1_lpi_1_dfm_3 <= _00638_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_uflow_2_lpi_1_dfm_3 <= 1'b0;
    else
      lut_lookup_lo_uflow_2_lpi_1_dfm_3 <= _00640_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_uflow_3_lpi_1_dfm_3 <= 1'b0;
    else
      lut_lookup_lo_uflow_3_lpi_1_dfm_3 <= _00642_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_uflow_lpi_1_dfm_3 <= 1'b0;
    else
      lut_lookup_lo_uflow_lpi_1_dfm_3 <= _00644_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2 <= 1'b0;
    else
      lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2 <= _00512_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_13 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_13 <= _00631_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_13 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_13 <= _00628_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lut_lookup_else_1_and_1_itm_2 <= 1'b0;
    else
      lut_lookup_else_1_lut_lookup_else_1_and_1_itm_2 <= _00468_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lut_lookup_else_1_and_4_itm_2 <= 1'b0;
    else
      lut_lookup_else_1_lut_lookup_else_1_and_4_itm_2 <= _00469_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2 <= 1'b0;
    else
      lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2 <= _00513_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2 <= 1'b0;
    else
      lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2 <= _00514_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2 <= 1'b0;
    else
      lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2 <= _00511_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_13 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_lpi_1_dfm_13 <= _00637_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_13 <= 8'b00000000;
    else
      lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_13 <= _00634_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lut_lookup_else_1_and_7_itm_2 <= 1'b0;
    else
      lut_lookup_else_1_lut_lookup_else_1_and_7_itm_2 <= _00470_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_1_lut_lookup_else_1_and_10_itm_2 <= 1'b0;
    else
      lut_lookup_else_1_lut_lookup_else_1_and_10_itm_2 <= _00467_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_uflow_1_lpi_1_dfm_6 <= 1'b0;
    else
      lut_lookup_le_uflow_1_lpi_1_dfm_6 <= _00618_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_uflow_2_lpi_1_dfm_6 <= 1'b0;
    else
      lut_lookup_le_uflow_2_lpi_1_dfm_6 <= _00619_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_uflow_3_lpi_1_dfm_6 <= 1'b0;
    else
      lut_lookup_le_uflow_3_lpi_1_dfm_6 <= _00620_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_uflow_lpi_1_dfm_6 <= 1'b0;
    else
      lut_lookup_le_uflow_lpi_1_dfm_6 <= _00621_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2 <= _00173_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_10_land_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_10_land_lpi_1_dfm_6 <= _00201_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 <= 1'b0;
    else
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 <= _00438_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_else_lo_fra_sva_4 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_if_1_else_lo_fra_sva_4 <= _00549_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_sva_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_sva_2 <= _00181_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_6_land_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_6_land_lpi_1_dfm_7 <= _00237_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 <= 1'b0;
    else
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 <= _00440_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_else_le_fra_sva_4 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_else_if_else_le_fra_sva_4 <= _00526_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_2_else_else_if_mux_26_itm_1 <= 1'b0;
    else
      lut_lookup_else_2_else_else_if_mux_26_itm_1 <= _00489_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_1_lpi_1_dfm_5 <= 1'b0;
    else
      lut_lookup_if_1_lor_1_lpi_1_dfm_5 <= _00551_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_7_lpi_1_dfm_5 <= 1'b0;
    else
      lut_lookup_if_1_lor_7_lpi_1_dfm_5 <= _00560_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2 <= _00172_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_10_land_3_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_10_land_3_lpi_1_dfm_6 <= _00199_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 <= 1'b0;
    else
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 <= _00412_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_else_lo_fra_3_sva_4 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_if_1_else_lo_fra_3_sva_4 <= _00548_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_1_lpi_1_dfm_6 <= 1'b0;
    else
      lut_lookup_else_if_lor_1_lpi_1_dfm_6 <= _00528_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_7_lpi_1_dfm_6 <= 1'b0;
    else
      lut_lookup_else_if_lor_7_lpi_1_dfm_6 <= _00537_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_3_sva_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_3_sva_2 <= _00180_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_6_land_3_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_6_land_3_lpi_1_dfm_7 <= _00235_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 <= 1'b0;
    else
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 <= _00414_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_else_le_fra_3_sva_4 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_else_if_else_le_fra_3_sva_4 <= _00525_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_2_else_else_if_mux_19_itm_1 <= 1'b0;
    else
      lut_lookup_else_2_else_else_if_mux_19_itm_1 <= _00488_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2 <= _00171_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_10_land_2_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_10_land_2_lpi_1_dfm_6 <= _00197_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 <= 1'b0;
    else
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 <= _00387_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_else_lo_fra_2_sva_4 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_if_1_else_lo_fra_2_sva_4 <= _00547_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_6_lpi_1_dfm_st_3 <= 1'b0;
    else
      lut_lookup_else_if_lor_6_lpi_1_dfm_st_3 <= _00535_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_6_lpi_1_dfm_6 <= 1'b0;
    else
      lut_lookup_else_if_lor_6_lpi_1_dfm_6 <= _00534_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_2_sva_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_2_sva_2 <= _00179_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_6_land_2_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_6_land_2_lpi_1_dfm_7 <= _00233_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 <= 1'b0;
    else
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 <= _00389_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_else_le_fra_2_sva_4 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_else_if_else_le_fra_2_sva_4 <= _00524_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_2_else_else_if_mux_12_itm_1 <= 1'b0;
    else
      lut_lookup_else_2_else_else_if_mux_12_itm_1 <= _00487_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_5_lpi_1_dfm_st_4 <= 1'b0;
    else
      lut_lookup_if_1_lor_5_lpi_1_dfm_st_4 <= _00555_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_6_lpi_1_dfm_st_4 <= 1'b0;
    else
      lut_lookup_if_1_lor_6_lpi_1_dfm_st_4 <= _00558_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_7_lpi_1_dfm_st_4 <= 1'b0;
    else
      lut_lookup_if_1_lor_7_lpi_1_dfm_st_4 <= _00561_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_1_lpi_1_dfm_st_4 <= 1'b0;
    else
      lut_lookup_if_1_lor_1_lpi_1_dfm_st_4 <= _00552_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_6_lpi_1_dfm_5 <= 1'b0;
    else
      lut_lookup_if_1_lor_6_lpi_1_dfm_5 <= _00557_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_lor_5_lpi_1_dfm_5 <= 1'b0;
    else
      lut_lookup_if_1_lor_5_lpi_1_dfm_5 <= _00554_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2 <= _00170_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_10_land_1_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_10_land_1_lpi_1_dfm_6 <= _00195_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 <= 1'b0;
    else
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2 <= _00362_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_1_else_lo_fra_1_sva_4 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_if_1_else_lo_fra_1_sva_4 <= _00546_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_precision_1_sva_st_72 <= 2'b00;
    else
      cfg_precision_1_sva_st_72 <= _00304_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_5_lpi_1_dfm_st_3 <= 1'b0;
    else
      lut_lookup_else_if_lor_5_lpi_1_dfm_st_3 <= _00532_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_7_lpi_1_dfm_st_3 <= 1'b0;
    else
      lut_lookup_else_if_lor_7_lpi_1_dfm_st_3 <= _00538_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_1_lpi_1_dfm_st_3 <= 1'b0;
    else
      lut_lookup_else_if_lor_1_lpi_1_dfm_st_3 <= _00529_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_lor_5_lpi_1_dfm_6 <= 1'b0;
    else
      lut_lookup_else_if_lor_5_lpi_1_dfm_6 <= _00531_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_1_sva_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_1_sva_2 <= _00178_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_6_land_1_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_6_land_1_lpi_1_dfm_7 <= _00231_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 <= 1'b0;
    else
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2 <= _00364_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_if_else_le_fra_1_sva_4 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_else_if_else_le_fra_1_sva_4 <= _00523_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_2_else_else_if_mux_5_itm_1 <= 1'b0;
    else
      lut_lookup_else_2_else_else_if_mux_5_itm_1 <= _00490_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_unequal_tmp_13 <= 1'b0;
    else
      lut_lookup_else_unequal_tmp_13 <= _00544_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_fraction_lpi_1_dfm_9 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_lo_fraction_lpi_1_dfm_9 <= _00625_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_lpi_1_dfm_26 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_lpi_1_dfm_26 <= _00614_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_lpi_1_dfm_21 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_le_fraction_lpi_1_dfm_21 <= _00596_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_lpi_1_dfm_28 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_lpi_1_dfm_28 <= _00616_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_lpi_1_dfm_22 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_le_fraction_lpi_1_dfm_22 <= _00597_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_lpi_1_dfm_29 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_lpi_1_dfm_29 <= _00617_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_fraction_3_lpi_1_dfm_9 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_lo_fraction_3_lpi_1_dfm_9 <= _00624_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_26 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_26 <= _00609_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_3_lpi_1_dfm_21 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_le_fraction_3_lpi_1_dfm_21 <= _00593_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_28 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_28 <= _00611_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_3_lpi_1_dfm_22 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_le_fraction_3_lpi_1_dfm_22 <= _00594_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_29 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_29 <= _00612_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_fraction_2_lpi_1_dfm_9 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_lo_fraction_2_lpi_1_dfm_9 <= _00623_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_26 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_26 <= _00604_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_2_lpi_1_dfm_21 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_le_fraction_2_lpi_1_dfm_21 <= _00590_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_28 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_28 <= _00606_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_2_lpi_1_dfm_22 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_le_fraction_2_lpi_1_dfm_22 <= _00591_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_29 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_29 <= _00607_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_fraction_1_lpi_1_dfm_9 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_lo_fraction_1_lpi_1_dfm_9 <= _00622_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_26 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_26 <= _00599_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_1_lpi_1_dfm_21 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_le_fraction_1_lpi_1_dfm_21 <= _00587_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_28 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_28 <= _00601_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_1_lpi_1_dfm_22 <= 35'b00000000000000000000000000000000000;
    else
      lut_lookup_le_fraction_1_lpi_1_dfm_22 <= _00588_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_29 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_29 <= _00602_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_function_1_sva_10 <= 1'b0;
    else
      cfg_lut_le_function_1_sva_10 <= _00271_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_uflow_priority_1_sva_10 <= 1'b0;
    else
      cfg_lut_uflow_priority_1_sva_10 <= _00295_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_oflow_priority_1_sva_10 <= 1'b0;
    else
      cfg_lut_oflow_priority_1_sva_10 <= _00290_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_hybrid_priority_1_sva_10 <= 1'b0;
    else
      cfg_lut_hybrid_priority_1_sva_10 <= _00266_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_in_data_sva_158 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      lut_in_data_sva_158 <= _00357_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_unequal_tmp_13 <= 1'b0;
    else
      lut_lookup_unequal_tmp_13 <= _00646_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_uflow_1_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_lo_uflow_1_lpi_1_dfm_4 <= _00639_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_and_svs_2 <= 1'b0;
    else
      lut_lookup_1_and_svs_2 <= _00369_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_uflow_2_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_lo_uflow_2_lpi_1_dfm_4 <= _00641_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_and_svs_2 <= 1'b0;
    else
      lut_lookup_2_and_svs_2 <= _00394_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_uflow_3_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_lo_uflow_3_lpi_1_dfm_4 <= _00643_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_and_svs_2 <= 1'b0;
    else
      lut_lookup_3_and_svs_2 <= _00419_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_lo_uflow_lpi_1_dfm_4 <= 1'b0;
    else
      lut_lookup_lo_uflow_lpi_1_dfm_4 <= _00645_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_and_svs_2 <= 1'b0;
    else
      lut_lookup_4_and_svs_2 <= _00445_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_precision_1_sva_st_107 <= 2'b00;
    else
      cfg_precision_1_sva_st_107 <= _00301_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_lpi_1_dfm_16_34_12_1 <= 23'b00000000000000000000000;
    else
      lut_lookup_le_fraction_lpi_1_dfm_16_34_12_1 <= _00595_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_3_lpi_1_dfm_16_34_12_1 <= 23'b00000000000000000000000;
    else
      lut_lookup_le_fraction_3_lpi_1_dfm_16_34_12_1 <= _00592_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_2_lpi_1_dfm_16_34_12_1 <= 23'b00000000000000000000000;
    else
      lut_lookup_le_fraction_2_lpi_1_dfm_16_34_12_1 <= _00589_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_fraction_1_lpi_1_dfm_16_34_12_1 <= 23'b00000000000000000000000;
    else
      lut_lookup_le_fraction_1_lpi_1_dfm_16_34_12_1 <= _00586_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_if_unequal_cse <= 1'b0;
    else
      reg_lut_lookup_if_unequal_cse <= _00727_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_5 <= 1'b0;
    else
      main_stage_v_5 <= _00651_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 <= 1'b0;
    else
      lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 <= _00449_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= 8'b00000000;
    else
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= _00437_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_4_itm_1_0_1 <= 1'b0;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_4_itm_1_0_1 <= _00168_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_sva_st_3 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_sva_st_3 <= _00502_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= 8'b00000000;
    else
      lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= _00439_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_4_itm_1_0_1 <= 1'b0;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_4_itm_1_0_1 <= _00176_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_sva_st_3 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_sva_st_3 <= _00581_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 <= 1'b0;
    else
      lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 <= _00452_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 <= 1'b0;
    else
      lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 <= _00423_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= 8'b00000000;
    else
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= _00411_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_3_itm_1_0_1 <= 1'b0;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_3_itm_1_0_1 <= _00167_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_3_sva_st_3 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_3_sva_st_3 <= _00499_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= 8'b00000000;
    else
      lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= _00413_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_3_itm_1_0_1 <= 1'b0;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_3_itm_1_0_1 <= _00175_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3 <= _00578_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 <= 1'b0;
    else
      lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 <= _00426_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 <= 1'b0;
    else
      lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 <= _00398_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= 8'b00000000;
    else
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= _00386_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_2_itm_1_0_1 <= 1'b0;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_2_itm_1_0_1 <= _00166_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_2_sva_st_3 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_2_sva_st_3 <= _00496_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= 8'b00000000;
    else
      lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= _00388_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_2_itm_1_0_1 <= 1'b0;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_2_itm_1_0_1 <= _00174_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3 <= _00575_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 <= 1'b0;
    else
      lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 <= _00401_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 <= 1'b0;
    else
      lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3 <= _00373_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= 8'b00000000;
    else
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 <= _00361_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_itm_1_0_1 <= 1'b0;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_itm_1_0_1 <= _00169_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_else_else_asn_mdf_1_sva_st_3 <= 1'b0;
    else
      lut_lookup_else_else_else_asn_mdf_1_sva_st_3 <= _00493_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= 8'b00000000;
    else
      lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2 <= _00363_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_1_0_1 <= 1'b0;
    else
      FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_1_0_1 <= _00177_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_else_unequal_tmp_18 <= 1'b0;
    else
      lut_lookup_else_unequal_tmp_18 <= _00545_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_lpi_1_dfm_25 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_lpi_1_dfm_25 <= _00613_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_lpi_1_dfm_27 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_lpi_1_dfm_27 <= _00615_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_25 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_25 <= _00608_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_27 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_3_lpi_1_dfm_27 <= _00610_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_25 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_25 <= _00603_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_27 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_2_lpi_1_dfm_27 <= _00605_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_25 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_25 <= _00598_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_27 <= 6'b000000;
    else
      lut_lookup_le_index_0_5_0_1_lpi_1_dfm_27 <= _00600_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_uflow_priority_1_sva_9 <= 1'b0;
    else
      cfg_lut_uflow_priority_1_sva_9 <= _00299_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_oflow_priority_1_sva_9 <= 1'b0;
    else
      cfg_lut_oflow_priority_1_sva_9 <= _00294_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_hybrid_priority_1_sva_9 <= 1'b0;
    else
      cfg_lut_hybrid_priority_1_sva_9 <= _00270_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_in_data_sva_157 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      lut_in_data_sva_157 <= _00356_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_precision_1_sva_st_71 <= 2'b00;
    else
      cfg_precision_1_sva_st_71 <= _00303_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_function_1_sva_st_42 <= 1'b0;
    else
      cfg_lut_le_function_1_sva_st_42 <= _00273_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_if_else_slc_32_svs_st_5 <= 1'b0;
    else
      lut_lookup_1_if_else_slc_32_svs_st_5 <= _00382_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_if_else_slc_32_svs_st_5 <= 1'b0;
    else
      lut_lookup_2_if_else_slc_32_svs_st_5 <= _00407_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_if_else_slc_32_svs_st_5 <= 1'b0;
    else
      lut_lookup_3_if_else_slc_32_svs_st_5 <= _00432_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_if_else_slc_32_svs_st_5 <= 1'b0;
    else
      lut_lookup_4_if_else_slc_32_svs_st_5 <= _00458_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3 <= _00572_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 <= 1'b0;
    else
      lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 <= _00376_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_index_offset_1_sva_7 <= 8'b00000000;
    else
      cfg_lut_le_index_offset_1_sva_7 <= _00277_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_4 <= 1'b0;
    else
      main_stage_v_4 <= _00650_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_61_itm_3 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_61_itm_3 <= _00149_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12 <= _00153_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_49U_24U_2_else_carry_sva_2 <= 1'b0;
    else
      FpMantRNE_49U_24U_2_else_carry_sva_2 <= _00189_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 <= 23'b00000000000000000000000;
    else
      lut_lookup_4_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 <= _00443_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_61_itm_4 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_61_itm_4 <= _00117_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm <= 6'b000000;
    else
      reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm <= _00658_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm <= 2'b00;
    else
      reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm <= _00659_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_49U_24U_1_else_carry_sva_2 <= 1'b0;
    else
      FpMantRNE_49U_24U_1_else_carry_sva_2 <= _00185_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 <= 23'b00000000000000000000000;
    else
      lut_lookup_4_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 <= _00441_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm <= 2'b00;
    else
      reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm <= _00725_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm <= 1'b0;
    else
      reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm <= _00726_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_lpi_1_dfm_8 <= _00212_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_45_itm_3 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_45_itm_3 <= _00146_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12 <= _00152_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_49U_24U_2_else_carry_3_sva_2 <= 1'b0;
    else
      FpMantRNE_49U_24U_2_else_carry_3_sva_2 <= _00188_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 <= 23'b00000000000000000000000;
    else
      lut_lookup_3_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 <= _00417_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_45_itm_4 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_45_itm_4 <= _00114_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm <= 6'b000000;
    else
      reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm <= _00656_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm <= 2'b00;
    else
      reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm <= _00657_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_49U_24U_1_else_carry_3_sva_2 <= 1'b0;
    else
      FpMantRNE_49U_24U_1_else_carry_3_sva_2 <= _00184_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 <= 23'b00000000000000000000000;
    else
      lut_lookup_3_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 <= _00415_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm <= 2'b00;
    else
      reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm <= _00714_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm <= 1'b0;
    else
      reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm <= _00715_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 <= _00209_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_29_itm_3 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_29_itm_3 <= _00143_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 <= _00259_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2 <= 1'b0;
    else
      lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2 <= _00391_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_7 <= _00244_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_6 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_6 <= _00246_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12 <= _00151_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_49U_24U_2_else_carry_2_sva_2 <= 1'b0;
    else
      FpMantRNE_49U_24U_2_else_carry_2_sva_2 <= _00187_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 <= 23'b00000000000000000000000;
    else
      lut_lookup_2_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 <= _00392_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 <= 1'b0;
    else
      FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 <= _00103_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 <= 1'b0;
    else
      FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 <= _00104_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 <= 1'b0;
    else
      FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 <= _00105_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_29_itm_4 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_29_itm_4 <= _00111_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm <= 6'b000000;
    else
      reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm <= _00654_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm <= 2'b00;
    else
      reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm <= _00655_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_49U_24U_1_else_carry_2_sva_2 <= 1'b0;
    else
      FpMantRNE_49U_24U_1_else_carry_2_sva_2 <= _00183_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 <= 23'b00000000000000000000000;
    else
      lut_lookup_2_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 <= _00390_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm <= 2'b00;
    else
      reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm <= _00703_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm <= 1'b0;
    else
      reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm <= _00704_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 <= _00207_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 <= 1'b0;
    else
      FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 <= _00134_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 <= 1'b0;
    else
      FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 <= _00135_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 <= 1'b0;
    else
      FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 <= _00136_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 <= 1'b0;
    else
      FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 <= _00137_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_mux_13_itm_3 <= 1'b0;
    else
      FpAdd_8U_23U_2_mux_13_itm_3 <= _00139_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_lo_start_1_sva_3_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      cfg_lut_lo_start_1_sva_3_30_0_1 <= _00288_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12 <= _00150_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_49U_24U_2_else_carry_1_sva_2 <= 1'b0;
    else
      FpMantRNE_49U_24U_2_else_carry_1_sva_2 <= _00186_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 <= 23'b00000000000000000000000;
    else
      lut_lookup_1_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2 <= _00367_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 <= 1'b0;
    else
      FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 <= _00102_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_8_land_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_8U_23U_8_land_lpi_1_dfm_5 <= _00263_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_8_land_3_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_8U_23U_8_land_3_lpi_1_dfm_5 <= _00261_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2 <= 1'b0;
    else
      lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2 <= _00366_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_7 <= _00239_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2 <= 1'b0;
    else
      lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2 <= _00416_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_7 <= _00248_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2 <= 1'b0;
    else
      lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2 <= _00442_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_lpi_1_dfm_7 <= _00253_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_6 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_6 <= _00242_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_6 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_6 <= _00251_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_lpi_1_dfm_st_6 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_lpi_1_dfm_st_6 <= _00254_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= 1'b0;
    else
      reg_lut_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= _00685_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= 1'b0;
    else
      reg_lut_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= _00696_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= 1'b0;
    else
      reg_lut_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= _00707_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= 1'b0;
    else
      reg_lut_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= _00718_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 <= _00213_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 <= _00215_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 <= 1'b0;
    else
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 <= _00218_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_3_land_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_3_land_lpi_1_dfm_6 <= _00220_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_st_6 <= 1'b0;
    else
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_st_6 <= _00214_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_6 <= 1'b0;
    else
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_6 <= _00217_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_st_6 <= 1'b0;
    else
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_st_6 <= _00219_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_3_land_lpi_1_dfm_st_6 <= 1'b0;
    else
      IsNaN_8U_23U_3_land_lpi_1_dfm_st_6 <= _00221_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_mux_13_itm_4 <= 1'b0;
    else
      FpAdd_8U_23U_1_mux_13_itm_4 <= _00107_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm <= 6'b000000;
    else
      reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm <= _00652_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm <= 2'b00;
    else
      reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm <= _00653_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpMantRNE_49U_24U_1_else_carry_1_sva_2 <= 1'b0;
    else
      FpMantRNE_49U_24U_1_else_carry_1_sva_2 <= _00182_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 <= 23'b00000000000000000000000;
    else
      lut_lookup_1_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2 <= _00365_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm <= 2'b00;
    else
      reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm <= _00692_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm <= 1'b0;
    else
      reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm <= _00693_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 <= _00204_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_if_else_slc_32_svs_7 <= 1'b0;
    else
      lut_lookup_4_if_else_slc_32_svs_7 <= _00456_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_if_else_slc_32_svs_7 <= 1'b0;
    else
      lut_lookup_3_if_else_slc_32_svs_7 <= _00430_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_if_else_slc_32_svs_7 <= 1'b0;
    else
      lut_lookup_2_if_else_slc_32_svs_7 <= _00405_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_if_else_slc_32_svs_7 <= 1'b0;
    else
      lut_lookup_1_if_else_slc_32_svs_7 <= _00380_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_sva_3 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_sva_3 <= _00579_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_3_sva_3 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_3_sva_3 <= _00576_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_2_sva_3 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_2_sva_3 <= _00573_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_if_else_else_slc_10_mdf_1_sva_3 <= 1'b0;
    else
      lut_lookup_if_else_else_slc_10_mdf_1_sva_3 <= _00570_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_index_offset_1_sva_6 <= 8'b00000000;
    else
      cfg_lut_le_index_offset_1_sva_6 <= _00276_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_index_select_1_sva_6 <= 8'b00000000;
    else
      cfg_lut_le_index_select_1_sva_6 <= _00280_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_lo_index_select_1_sva_6 <= 8'b00000000;
    else
      cfg_lut_lo_index_select_1_sva_6 <= _00286_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_uflow_priority_1_sva_8 <= 1'b0;
    else
      cfg_lut_uflow_priority_1_sva_8 <= _00298_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_oflow_priority_1_sva_8 <= 1'b0;
    else
      cfg_lut_oflow_priority_1_sva_8 <= _00293_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_hybrid_priority_1_sva_8 <= 1'b0;
    else
      cfg_lut_hybrid_priority_1_sva_8 <= _00269_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_in_data_sva_156 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      lut_in_data_sva_156 <= _00355_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_precision_1_sva_st_70 <= 2'b00;
    else
      cfg_precision_1_sva_st_70 <= _00302_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_function_1_sva_st_41 <= 1'b0;
    else
      cfg_lut_le_function_1_sva_st_41 <= _00272_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_start_1_sva_3_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      cfg_lut_le_start_1_sva_3_30_0_1 <= _00282_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_3 <= 1'b0;
    else
      main_stage_v_3 <= _00649_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_int_mant_p1_sva_3 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_2_int_mant_p1_sva_3 <= _00129_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_int_mant_p1_sva_3 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_1_int_mant_p1_sva_3 <= _00097_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm <= 6'b000000;
    else
      reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm <= _00666_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_int_mant_p1_3_sva_3 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_2_int_mant_p1_3_sva_3 <= _00128_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_8_land_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_8U_23U_8_land_lpi_1_dfm_4 <= _00262_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 <= 1'b0;
    else
      IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 <= _00260_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5 <= _00163_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_qr_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_qr_lpi_1_dfm_5 <= _00165_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5 <= _00250_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse <= 1'b0;
    else
      reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse <= _00677_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_int_mant_p1_3_sva_3 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_1_int_mant_p1_3_sva_3 <= _00096_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm <= 6'b000000;
    else
      reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm <= _00664_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_int_mant_p1_2_sva_3 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_2_int_mant_p1_2_sva_3 <= _00127_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5 <= _00161_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5 <= _00245_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_int_mant_p1_2_sva_3 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_1_int_mant_p1_2_sva_3 <= _00095_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm <= 6'b000000;
    else
      reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm <= _00662_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm <= 2'b00;
    else
      reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm <= _00663_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm <= 2'b00;
    else
      reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm <= _00665_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm <= 2'b00;
    else
      reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm <= _00667_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_int_mant_p1_1_sva_3 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_2_int_mant_p1_1_sva_3 <= _00126_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_8_land_1_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_8_land_1_lpi_1_dfm_6 <= _00257_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5 <= _00159_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5 <= _00241_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_int_mant_p1_1_sva_3 <= 50'b00000000000000000000000000000000000000000000000000;
    else
      FpAdd_8U_23U_1_int_mant_p1_1_sva_3 <= _00094_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm <= 6'b000000;
    else
      reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm <= _00660_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm <= 2'b00;
    else
      reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm <= _00661_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_if_else_slc_32_svs_6 <= 1'b0;
    else
      lut_lookup_4_if_else_slc_32_svs_6 <= _00455_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_if_else_slc_32_svs_6 <= 1'b0;
    else
      lut_lookup_3_if_else_slc_32_svs_6 <= _00429_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_if_else_slc_32_svs_6 <= 1'b0;
    else
      lut_lookup_2_if_else_slc_32_svs_6 <= _00404_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_if_else_slc_32_svs_6 <= 1'b0;
    else
      lut_lookup_1_if_else_slc_32_svs_6 <= _00379_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_index_offset_1_sva_5 <= 8'b00000000;
    else
      cfg_lut_le_index_offset_1_sva_5 <= _00275_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_index_select_1_sva_5 <= 8'b00000000;
    else
      cfg_lut_le_index_select_1_sva_5 <= _00279_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_lo_index_select_1_sva_5 <= 8'b00000000;
    else
      cfg_lut_lo_index_select_1_sva_5 <= _00285_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_uflow_priority_1_sva_7 <= 1'b0;
    else
      cfg_lut_uflow_priority_1_sva_7 <= _00297_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_oflow_priority_1_sva_7 <= 1'b0;
    else
      cfg_lut_oflow_priority_1_sva_7 <= _00292_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_hybrid_priority_1_sva_7 <= 1'b0;
    else
      cfg_lut_hybrid_priority_1_sva_7 <= _00268_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_in_data_sva_155 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      lut_in_data_sva_155 <= _00354_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_start_1_sva_2_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      cfg_lut_le_start_1_sva_2_30_0_1 <= _00281_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_lo_start_1_sva_2_30_0_1 <= 31'b0000000000000000000000000000000;
    else
      cfg_lut_lo_start_1_sva_2_30_0_1 <= _00287_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_cfg_precision_1_sva_st_13_cse_1 <= 2'b00;
    else
      reg_cfg_precision_1_sva_st_13_cse_1 <= _00681_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_cfg_lut_le_function_1_sva_st_20_cse <= 1'b0;
    else
      reg_cfg_lut_le_function_1_sva_st_20_cse <= _00679_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_2 <= 1'b0;
    else
      main_stage_v_2 <= _00648_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_8_land_2_lpi_1_dfm_5 <= 1'b0;
    else
      IsNaN_8U_23U_8_land_2_lpi_1_dfm_5 <= _00258_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 <= 1'b0;
    else
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_6 <= _00205_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_a_right_shift_qr_sva_3 <= 8'b00000000;
    else
      FpAdd_8U_23U_1_a_right_shift_qr_sva_3 <= _00093_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_a_right_shift_qr_3_sva_3 <= 8'b00000000;
    else
      FpAdd_8U_23U_1_a_right_shift_qr_3_sva_3 <= _00092_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_a_right_shift_qr_2_sva_3 <= 8'b00000000;
    else
      FpAdd_8U_23U_1_a_right_shift_qr_2_sva_3 <= _00091_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_qr_3_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_1_qr_3_lpi_1_dfm_5 <= _00119_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_qr_4_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_1_qr_4_lpi_1_dfm_5 <= _00120_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_1_qr_lpi_1_dfm_5 <= 8'b00000000;
    else
      FpAdd_8U_23U_1_qr_lpi_1_dfm_5 <= _00121_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= 1'b0;
    else
      lut_lookup_2_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= _00385_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4 <= 1'b0;
    else
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4 <= _00216_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4 <= _00249_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_2_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse <= 1'b0;
    else
      reg_lut_lookup_2_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse <= _00695_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse <= 1'b0;
    else
      reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse <= _00694_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse <= 1'b0;
    else
      reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse <= _00705_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse <= 1'b0;
    else
      reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse <= _00706_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse <= 1'b0;
    else
      reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse <= _00716_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse <= 1'b0;
    else
      reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse <= _00717_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse <= 1'b0;
    else
      reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse <= _00676_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_a_right_shift_qr_1_sva_3 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_a_right_shift_qr_1_sva_3 <= _00122_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      FpAdd_8U_23U_2_qr_2_lpi_1_dfm_4 <= 8'b00000000;
    else
      FpAdd_8U_23U_2_qr_2_lpi_1_dfm_4 <= _00158_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= 1'b0;
    else
      lut_lookup_1_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2 <= _00360_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4 <= 1'b0;
    else
      IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4 <= _00240_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_1_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse <= 1'b0;
    else
      reg_lut_lookup_1_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse <= _00684_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse <= 1'b0;
    else
      reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse <= _00683_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_4_if_else_slc_32_svs_5 <= 1'b0;
    else
      lut_lookup_4_if_else_slc_32_svs_5 <= _00454_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_3_if_else_slc_32_svs_5 <= 1'b0;
    else
      lut_lookup_3_if_else_slc_32_svs_5 <= _00428_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_2_if_else_slc_32_svs_5 <= 1'b0;
    else
      lut_lookup_2_if_else_slc_32_svs_5 <= _00403_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_lookup_1_if_else_slc_32_svs_5 <= 1'b0;
    else
      lut_lookup_1_if_else_slc_32_svs_5 <= _00378_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_start_1_sva_41 <= 32'd0;
    else
      cfg_lut_le_start_1_sva_41 <= _00283_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_lo_start_1_sva_41 <= 32'd0;
    else
      cfg_lut_lo_start_1_sva_41 <= _00289_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_index_offset_1_sva_4 <= 8'b00000000;
    else
      cfg_lut_le_index_offset_1_sva_4 <= _00274_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_le_index_select_1_sva_4 <= 8'b00000000;
    else
      cfg_lut_le_index_select_1_sva_4 <= _00278_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_lo_index_select_1_sva_4 <= 8'b00000000;
    else
      cfg_lut_lo_index_select_1_sva_4 <= _00284_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_uflow_priority_1_sva_6 <= 1'b0;
    else
      cfg_lut_uflow_priority_1_sva_6 <= _00296_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_oflow_priority_1_sva_6 <= 1'b0;
    else
      cfg_lut_oflow_priority_1_sva_6 <= _00291_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cfg_lut_hybrid_priority_1_sva_6 <= 1'b0;
    else
      cfg_lut_hybrid_priority_1_sva_6 <= _00267_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      lut_in_data_sva_154 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      lut_in_data_sva_154 <= _00353_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_cfg_precision_1_sva_st_12_cse_1 <= 2'b00;
    else
      reg_cfg_precision_1_sva_st_12_cse_1 <= _00680_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_cfg_lut_le_function_1_sva_st_19_cse <= 1'b0;
    else
      reg_cfg_lut_le_function_1_sva_st_19_cse <= _00678_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      main_stage_v_1 <= 1'b0;
    else
      main_stage_v_1 <= _00647_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg_chn_lut_out_rsci_ld_core_psct_cse <= 1'b0;
    else
      reg_chn_lut_out_rsci_ld_core_psct_cse <= _00682_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_315 <= 1'b0;
    else
      chn_lut_out_rsci_d_315 <= _00339_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_314 <= 1'b0;
    else
      chn_lut_out_rsci_d_314 <= _00338_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_313 <= 1'b0;
    else
      chn_lut_out_rsci_d_313 <= _00337_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_279 <= 1'b0;
    else
      chn_lut_out_rsci_d_279 <= _00323_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_275 <= 1'b0;
    else
      chn_lut_out_rsci_d_275 <= _00319_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_306 <= 1'b0;
    else
      chn_lut_out_rsci_d_306 <= _00335_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_305 <= 1'b0;
    else
      chn_lut_out_rsci_d_305 <= _00334_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_304 <= 1'b0;
    else
      chn_lut_out_rsci_d_304 <= _00333_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_278 <= 1'b0;
    else
      chn_lut_out_rsci_d_278 <= _00322_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_274 <= 1'b0;
    else
      chn_lut_out_rsci_d_274 <= _00318_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_297 <= 1'b0;
    else
      chn_lut_out_rsci_d_297 <= _00331_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_296 <= 1'b0;
    else
      chn_lut_out_rsci_d_296 <= _00330_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_295 <= 1'b0;
    else
      chn_lut_out_rsci_d_295 <= _00329_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_277 <= 1'b0;
    else
      chn_lut_out_rsci_d_277 <= _00321_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_273 <= 1'b0;
    else
      chn_lut_out_rsci_d_273 <= _00317_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_288 <= 1'b0;
    else
      chn_lut_out_rsci_d_288 <= _00327_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_287 <= 1'b0;
    else
      chn_lut_out_rsci_d_287 <= _00326_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_286 <= 1'b0;
    else
      chn_lut_out_rsci_d_286 <= _00325_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_276 <= 1'b0;
    else
      chn_lut_out_rsci_d_276 <= _00320_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_272 <= 1'b0;
    else
      chn_lut_out_rsci_d_272 <= _00316_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_323 <= 1'b0;
    else
      chn_lut_out_rsci_d_323 <= _00347_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_322 <= 1'b0;
    else
      chn_lut_out_rsci_d_322 <= _00346_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_321 <= 1'b0;
    else
      chn_lut_out_rsci_d_321 <= _00345_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_320 <= 1'b0;
    else
      chn_lut_out_rsci_d_320 <= _00344_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_319 <= 1'b0;
    else
      chn_lut_out_rsci_d_319 <= _00343_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_318 <= 1'b0;
    else
      chn_lut_out_rsci_d_318 <= _00342_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_317 <= 1'b0;
    else
      chn_lut_out_rsci_d_317 <= _00341_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_316 <= 1'b0;
    else
      chn_lut_out_rsci_d_316 <= _00340_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_312_307 <= 6'b000000;
    else
      chn_lut_out_rsci_d_312_307 <= _00336_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_303_298 <= 6'b000000;
    else
      chn_lut_out_rsci_d_303_298 <= _00332_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_294_289 <= 6'b000000;
    else
      chn_lut_out_rsci_d_294_289 <= _00328_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_285_280 <= 6'b000000;
    else
      chn_lut_out_rsci_d_285_280 <= _00324_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_271 <= 1'b0;
    else
      chn_lut_out_rsci_d_271 <= _00315_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_270 <= 1'b0;
    else
      chn_lut_out_rsci_d_270 <= _00314_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_269 <= 1'b0;
    else
      chn_lut_out_rsci_d_269 <= _00313_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_268 <= 1'b0;
    else
      chn_lut_out_rsci_d_268 <= _00312_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_267_140 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      chn_lut_out_rsci_d_267_140 <= _00311_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_139_117 <= 23'b00000000000000000000000;
    else
      chn_lut_out_rsci_d_139_117 <= _00310_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_116_105 <= 12'b000000000000;
    else
      chn_lut_out_rsci_d_116_105 <= _00308_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_104_82 <= 23'b00000000000000000000000;
    else
      chn_lut_out_rsci_d_104_82 <= _00307_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_81_70 <= 12'b000000000000;
    else
      chn_lut_out_rsci_d_81_70 <= _00351_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_69_47 <= 23'b00000000000000000000000;
    else
      chn_lut_out_rsci_d_69_47 <= _00350_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_46_35 <= 12'b000000000000;
    else
      chn_lut_out_rsci_d_46_35 <= _00349_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_34_12 <= 23'b00000000000000000000000;
    else
      chn_lut_out_rsci_d_34_12 <= _00348_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_d_11_0 <= 12'b000000000000;
    else
      chn_lut_out_rsci_d_11_0 <= _00309_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_in_rsci_ld_core_psct <= 1'b0;
    else
      chn_lut_in_rsci_ld_core_psct <= _00306_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_out_rsci_iswt0 <= 1'b0;
    else
      chn_lut_out_rsci_iswt0 <= _00352_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      chn_lut_in_rsci_iswt0 <= 1'b0;
    else
      chn_lut_in_rsci_iswt0 <= _00305_;
  assign z_out_3 = lut_lookup_else_2_if_mux_34_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_if_mux_34_nl = lut_lookup_else_2_else_else_else_and_7_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_le_miss_sva : cfg_lut_oflow_priority_1_sva_10;
  assign mux_1297_nl = lut_lookup_else_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_201 : mux_1298_nl;
  assign mux_1298_nl = cfg_lut_le_function_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_882_nl : and_tmp_201;
  assign z_out_2 = lut_lookup_else_2_if_mux_33_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_if_mux_33_nl = lut_lookup_else_2_else_else_else_and_6_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_le_miss_3_sva : cfg_lut_oflow_priority_1_sva_10;
  assign mux_1294_nl = cfg_lut_le_function_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1295_nl : nand_118_nl;
  assign mux_1295_nl = lut_lookup_else_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nand_117_nl : or_2090_nl;
  assign z_out_1 = lut_lookup_else_2_if_mux_32_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_if_mux_32_nl = lut_lookup_else_2_else_else_else_and_5_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_le_miss_2_sva : cfg_lut_oflow_priority_1_sva_10;
  assign mux_1291_nl = cfg_lut_le_function_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1292_nl : nand_116_nl;
  assign mux_1292_nl = lut_lookup_else_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nand_115_nl : or_2089_nl;
  assign z_out = lut_lookup_else_2_if_mux_31_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_if_mux_31_nl = lut_lookup_else_2_else_else_else_and_4_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_le_miss_1_sva : cfg_lut_oflow_priority_1_sva_10;
  assign mux_1288_nl = cfg_lut_le_function_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1289_nl : nand_114_nl;
  assign mux_1289_nl = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nand_113_nl : or_2088_nl;
  assign mux_1118_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_178 : mux_tmp_1101;
  assign mux_1112_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_1104 : mux_982_cse;
  assign mux_1110_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_448_nl : nor_449_nl;
  assign mux_1107_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_450_nl : and_773_nl;
  assign mux_1104_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_451_nl : and_774_nl;
  assign mux_1103_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_1101 : and_42_cse;
  assign mux_1101_nl = or_1460_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1450 : mux_1100_nl;
  assign mux_1100_nl = FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1099_nl : or_tmp_1450;
  assign mux_1099_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nand_33_nl : or_1830_nl;
  assign mux_1098_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1458_nl : or_tmp_1250;
  assign mux_1097_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_236_nl : and_tmp_124;
  assign mux_1096_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1094_nl : mux_1095_nl;
  assign mux_1095_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_235_nl : nor_454_nl;
  assign mux_1094_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_233_nl : nor_453_nl;
  assign lut_lookup_else_else_else_lut_lookup_else_else_else_and_7_nl = lut_lookup_4_else_else_else_if_acc_nl[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_sva[5:0] : 6'b000000;
  assign mux_1093_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1450_nl : or_tmp_1181;
  assign mux_1092_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_232_nl : and_tmp_113;
  assign mux_1091_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1088_nl : mux_1090_nl;
  assign mux_1090_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_230_nl : nor_564_cse;
  assign mux_1088_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_228_nl : nor_455_nl;
  assign lut_lookup_else_else_else_lut_lookup_else_else_else_and_5_nl = lut_lookup_3_else_else_else_if_acc_nl[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_3_sva[5:0] : 6'b000000;
  assign mux_1086_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1440_nl : nand_tmp_22;
  assign mux_1085_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_226_nl : and_tmp_103;
  assign mux_1084_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1081_nl : mux_1083_nl;
  assign mux_1083_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_224_nl : nor_588_cse;
  assign mux_1081_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_222_nl : nor_459_nl;
  assign lut_lookup_else_else_else_lut_lookup_else_else_else_and_3_nl = lut_lookup_2_else_else_else_if_acc_nl[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_2_sva[5:0] : 6'b000000;
  assign mux_1079_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1431_nl : or_tmp_1043;
  assign mux_1078_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_221_nl : and_tmp_92;
  assign mux_1077_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1075_nl : mux_1076_nl;
  assign mux_1076_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_220_nl : nor_464_nl;
  assign mux_1075_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_219_nl : nor_463_nl;
  assign lut_lookup_else_else_else_lut_lookup_else_else_else_and_1_nl = lut_lookup_1_else_else_else_if_acc_nl[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_1_sva[5:0] : 6'b000000;
  assign mux_1073_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_467_nl : nor_468_nl;
  assign mux_1071_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_470_nl : nor_471_nl;
  assign mux_1070_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_472_nl : nor_473_nl;
  assign mux_1069_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_475_nl : mux_1068_nl;
  assign mux_1068_nl = reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_476_nl : nor_477_nl;
  assign mux_1066_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_480_nl : nor_481_nl;
  assign mux_1064_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_483_nl : nor_484_nl;
  assign mux_1063_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_485_nl : nor_486_nl;
  assign mux_1062_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_487_nl : nor_488_nl;
  assign mux_1061_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_489_nl : nor_490_nl;
  assign mux_1060_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_491_nl : nor_492_nl;
  assign mux_1059_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_493_nl : nor_494_nl;
  assign mux_1058_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_495_nl : mux_1057_nl;
  assign mux_1057_nl = IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_496_nl : nor_497_nl;
  assign mux_1055_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_42_cse : mux_793_cse;
  assign mux_1051_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_982_cse : and_tmp_6;
  assign mux_1049_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1146_nl : mux_959_cse;
  assign mux_nl = or_66_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : and_215_nl;
  assign mux_1033_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_500_nl : mux_1032_nl;
  assign mux_1032_nl = _03087_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_503_nl : nor_501_nl;
  assign mux_1031_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1148_nl : mux_900_cse;
  assign mux_1267_nl = or_66_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : and_204_nl;
  assign mux_1015_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_506_nl : mux_1014_nl;
  assign mux_1014_nl = _03081_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_509_nl : nor_507_nl;
  assign mux_1013_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1149_nl : mux_845_cse;
  assign mux_1268_nl = or_66_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : and_193_nl;
  assign mux_997_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_512_nl : mux_996_nl;
  assign mux_996_nl = _03075_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_515_nl : nor_513_nl;
  assign mux_995_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1147_nl : mux_789_cse;
  assign mux_1266_nl = or_66_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : and_179_nl;
  assign mux_986_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_178_cse : mux_851_cse;
  assign mux_981_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_518_nl : mux_980_nl;
  assign mux_980_nl = _03069_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_521_nl : nor_519_nl;
  assign mux_975_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_130 : and_tmp_131;
  assign mux_1252_nl = or_2035_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_825_nl : nand_nl;
  assign mux_971_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1250 : or_1252_nl;
  assign mux_969_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_427 : or_tmp_623;
  assign mux_962_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_959_cse : mux_961_nl;
  assign mux_961_nl = and_811_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : and_166_nl;
  assign mux_949_nl = cfg_precision_1_sva_st_71[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : nor_526_cse;
  assign mux_955_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_124 : and_163_nl;
  assign mux_954_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_528_nl : nor_529_nl;
  assign mux_953_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_771_cse : and_1174_nl;
  assign mux_1283_nl = or_2087_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : nor_526_cse;
  assign mux_945_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1151_nl : mux_944_nl;
  assign mux_944_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_612_cse : mux_943_nl;
  assign mux_943_nl = and_804_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_755_cse : _00027_;
  assign mux_1270_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : and_160_nl;
  assign mux_936_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1153_nl : _00031_;
  assign mux_935_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_978_cse : mux_934_nl;
  assign mux_934_nl = or_1213_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_993 : mux_933_nl;
  assign mux_933_nl = lut_lookup_4_if_else_slc_32_svs_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00025_ : or_tmp_993;
  assign mux_1271_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : nor_540_nl;
  assign mux_926_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00030_ : and_1176_nl;
  assign mux_1284_nl = or_1202_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_544_nl : main_stage_v_4;
  assign mux_916_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_158_nl : and_tmp_119;
  assign mux_1251_nl = or_2025_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_827_nl : nand_102_nl;
  assign mux_912_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1181 : or_1183_nl;
  assign mux_910_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_395 : or_tmp_573;
  assign mux_903_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_900_cse : mux_902_nl;
  assign mux_902_nl = and_811_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : mux_901_nl;
  assign mux_901_nl = cfg_precision_1_sva_st_71[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_281 : nor_549_nl;
  assign mux_896_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_113 : and_152_nl;
  assign mux_895_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_551_nl : nor_552_nl;
  assign mux_887_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1156_nl : mux_886_nl;
  assign mux_886_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_612_cse : mux_885_nl;
  assign mux_885_nl = and_808_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_755_cse : _00027_;
  assign mux_880_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : and_149_nl;
  assign mux_878_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1158_nl : _00029_;
  assign mux_877_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_978_cse : mux_876_nl;
  assign mux_876_nl = or_1142_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_993 : mux_875_nl;
  assign mux_875_nl = lut_lookup_3_if_else_slc_32_svs_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00025_ : or_tmp_993;
  assign mux_870_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : nor_564_cse;
  assign mux_861_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_6 : mux_805_cse;
  assign mux_859_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_147_nl : and_tmp_108;
  assign mux_1250_nl = _03700_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1249_nl : or_tmp_1720;
  assign mux_1249_nl = and_1140_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1720 : and_1089_nl;
  assign mux_855_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nand_tmp_22 : or_1113_nl;
  assign mux_854_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_363 : mux_tmp_301;
  assign mux_848_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_845_cse : mux_847_nl;
  assign mux_847_nl = and_811_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : mux_846_nl;
  assign mux_846_nl = cfg_precision_1_sva_st_71[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_260 : nor_573_nl;
  assign mux_841_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_103 : and_142_nl;
  assign mux_840_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_575_nl : nor_576_nl;
  assign mux_832_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1160_nl : mux_831_nl;
  assign mux_831_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_612_cse : mux_830_nl;
  assign mux_830_nl = and_812_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_755_cse : _00027_;
  assign mux_825_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : and_138_nl;
  assign mux_823_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1162_nl : _00028_;
  assign mux_822_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_978_cse : mux_821_nl;
  assign mux_821_nl = or_1072_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_993 : mux_820_nl;
  assign mux_820_nl = lut_lookup_2_if_else_slc_32_svs_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00025_ : or_tmp_993;
  assign mux_815_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : nor_588_cse;
  assign mux_806_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_793_cse : mux_805_cse;
  assign mux_803_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_97 : and_tmp_98;
  assign mux_1248_nl = or_2007_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_2009_nl : mux_1247_nl;
  assign mux_1247_nl = cfg_precision_1_sva_st_70[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1716 : nor_830_nl;
  assign mux_799_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1043 : or_1045_nl;
  assign mux_798_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_331 : mux_tmp_279;
  assign mux_797_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_851_cse : mux_796_nl;
  assign mux_796_nl = and_814_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : and_134_cse;
  assign mux_792_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_789_cse : mux_791_nl;
  assign mux_791_nl = and_814_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : mux_790_nl;
  assign mux_790_nl = cfg_precision_1_sva_st_71[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_238 : nor_595_nl;
  assign mux_785_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_92 : and_131_nl;
  assign mux_784_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_815_nl : and_816_nl;
  assign mux_783_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_597_nl : nor_598_nl;
  assign mux_1246_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_833_nl : nor_831_nl;
  assign mux_1245_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1142_cse : nor_832_cse;
  assign mux_768_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1164_nl : mux_767_nl;
  assign mux_767_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_612_cse : mux_766_nl;
  assign mux_766_nl = and_819_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_755_cse : _00027_;
  assign mux_761_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : and_127_nl;
  assign mux_759_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_1166_nl : _00026_;
  assign mux_758_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_978_cse : mux_757_nl;
  assign mux_757_nl = or_990_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_993 : mux_756_nl;
  assign mux_756_nl = lut_lookup_1_if_else_slc_32_svs_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00025_ : or_tmp_993;
  assign mux_751_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : nor_616_nl;
  assign mux_739_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_737_nl : mux_738_nl;
  assign mux_738_nl = lut_lookup_if_1_lor_5_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_83 : main_stage_v_4;
  assign mux_737_nl = or_969_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_6 : main_stage_v_3;
  assign mux_732_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_730_nl : mux_731_nl;
  assign mux_731_nl = lut_lookup_if_1_lor_6_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_83 : main_stage_v_4;
  assign mux_730_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : nor_619_nl;
  assign mux_722_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_822_nl : mux_721_nl;
  assign mux_721_nl = lut_lookup_if_1_lor_7_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_83 : main_stage_v_4;
  assign mux_711_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_823_nl : mux_710_nl;
  assign mux_710_nl = lut_lookup_if_1_lor_1_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_83 : main_stage_v_4;
  assign mux_704_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_670_cse : mux_tmp_270;
  assign mux_700_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_118_nl : and_119_nl;
  assign mux_699_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_697_nl : _00024_;
  assign mux_698_nl = or_939_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_314 : nor_626_nl;
  assign mux_697_nl = lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_314 : nand_20_nl;
  assign mux_696_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_931_nl : _00023_;
  assign mux_695_nl = or_932_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1857_cse : nor_623_nl;
  assign mux_689_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_116_nl : and_117_nl;
  assign mux_688_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_686_nl : _00022_;
  assign mux_687_nl = or_923_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_314 : nor_631_nl;
  assign mux_686_nl = lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_314 : nand_19_nl;
  assign mux_685_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_915_nl : _00021_;
  assign mux_684_nl = or_916_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1857_cse : nor_628_nl;
  assign mux_678_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_114_nl : and_115_nl;
  assign mux_677_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_675_nl : _00020_;
  assign mux_676_nl = or_907_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_314 : nor_636_nl;
  assign mux_675_nl = lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_314 : nand_18_nl;
  assign mux_674_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_899_nl : _00019_;
  assign mux_673_nl = or_900_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1857_cse : nor_633_nl;
  assign mux_672_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_826_cse : main_stage_v_4;
  assign mux_667_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_112_nl : and_113_nl;
  assign mux_666_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_664_nl : _00018_;
  assign mux_665_nl = or_888_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_314 : nor_640_nl;
  assign mux_664_nl = lut_lookup_else_if_lor_1_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_885_nl : or_887_nl;
  assign mux_663_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_879_nl : _00017_;
  assign mux_662_nl = or_880_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1857_cse : nor_638_nl;
  assign mux_661_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_110_nl : and_111_nl;
  assign mux_660_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_108_nl : and_109_nl;
  assign mux_659_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_106_nl : and_tmp_69;
  assign mux_658_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_104_nl : and_105_nl;
  assign mux_657_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_102_nl : and_103_nl;
  assign mux_655_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_100_nl : and_101_nl;
  assign mux_654_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_98_nl : and_tmp_61;
  assign mux_548_nl = reg_cfg_precision_1_sva_st_12_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_1 : not_tmp_422;
  assign mux_653_nl = and_827_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_652_nl : nor_642_nl;
  assign mux_652_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_1 : and_tmp_59;
  assign mux_651_nl = _03413_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_650_nl : mux_645_nl;
  assign mux_650_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_649_nl : mux_tmp_643;
  assign mux_649_nl = or_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_647_nl : mux_646_nl;
  assign mux_647_nl = or_849_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : not_tmp_418;
  assign mux_646_nl = reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1688_cse : nand_17_nl;
  assign mux_534_nl = reg_cfg_precision_1_sva_st_12_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : not_tmp_418;
  assign mux_645_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_638_nl : mux_tmp_643;
  assign mux_638_nl = or_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_636_nl : mux_635_nl;
  assign mux_636_nl = or_849_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00003_ : not_tmp_412;
  assign mux_635_nl = reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1688_cse : nand_16_nl;
  assign mux_518_nl = reg_cfg_precision_1_sva_st_12_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : _00016_;
  assign mux_634_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_627_nl : mux_631_nl;
  assign mux_631_nl = or_1688_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : mux_628_nl;
  assign mux_628_nl = or_850_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : _00000_;
  assign mux_627_nl = or_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_625_nl : mux_624_nl;
  assign mux_625_nl = or_849_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_475 : not_tmp_394;
  assign mux_624_nl = IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1688_cse : nand_15_nl;
  assign mux_477_nl = reg_cfg_precision_1_sva_st_12_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_475 : not_tmp_394;
  assign mux_622_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_621_nl : mux_tmp_617;
  assign mux_621_nl = reg_cfg_precision_1_sva_st_12_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_618 : mux_620_nl;
  assign mux_620_nl = reg_cfg_precision_1_sva_st_12_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00015_ : mux_tmp_618;
  assign mux_611_nl = main_stage_v_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_839_nl : or_cse;
  assign mux_606_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_600_nl : mux_605_nl;
  assign mux_605_nl = or_26_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : mux_602_nl;
  assign mux_602_nl = main_stage_v_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_601_nl : or_1689_cse;
  assign mux_601_nl = or_829_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : _00000_;
  assign mux_600_nl = reg_cfg_precision_1_sva_st_12_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_596 : mux_599_nl;
  assign mux_599_nl = reg_cfg_precision_1_sva_st_12_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00014_ : mux_tmp_596;
  assign mux_598_nl = or_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_827_nl : main_stage_v_1;
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_9_nl = FpAdd_8U_23U_2_b_right_shift_qif_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) _00041_ : _00045_;
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_8_nl = FpAdd_8U_23U_2_b_right_shift_qif_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) chn_lut_in_rsci_d_mxwt[126:119] : cfg_lut_lo_start_rsci_d[30:23];
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_13_nl = FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) _00041_ : _00044_;
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_12_nl = FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) chn_lut_in_rsci_d_mxwt[94:87] : cfg_lut_lo_start_rsci_d[30:23];
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_15_nl = FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) _00041_ : _00042_;
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_14_nl = FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) chn_lut_in_rsci_d_mxwt[62:55] : cfg_lut_lo_start_rsci_d[30:23];
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_9_nl = FpAdd_8U_23U_b_right_shift_qif_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) _00043_ : _00040_;
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_8_nl = FpAdd_8U_23U_b_right_shift_qif_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) chn_lut_in_rsci_d_mxwt[30:23] : cfg_lut_le_start_rsci_d[30:23];
  assign mux_372_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_830_nl : mux_371_nl;
  assign mux_371_nl = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_5 : not_tmp_334;
  assign mux_349_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_623 : or_625_nl;
  assign mux_346_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_428 : or_620_nl;
  assign mux_344_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_428 : or_617_nl;
  assign mux_343_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_658_nl : nor_659_nl;
  assign mux_335_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_660_nl : nor_661_nl;
  assign mux_334_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_596_nl : or_tmp_598;
  assign mux_333_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_662_nl : nor_663_nl;
  assign mux_332_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_664_nl : nor_665_nl;
  assign mux_1178_nl = cfg_lut_hybrid_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1177_nl : and_459_nl;
  assign mux_1177_nl = cfg_lut_uflow_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1545 : _00013_;
  assign mux_325_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_573 : or_575_nl;
  assign mux_322_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_397 : or_569_nl;
  assign mux_320_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_397 : or_566_nl;
  assign mux_319_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_666_nl : nor_667_nl;
  assign mux_311_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_668_nl : nor_669_nl;
  assign mux_310_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_545_nl : or_tmp_547;
  assign mux_309_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_670_nl : nor_671_nl;
  assign mux_308_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_672_nl : nor_673_nl;
  assign mux_1165_nl = cfg_lut_hybrid_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1164_nl : and_455_nl;
  assign mux_1164_nl = cfg_lut_uflow_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1534 : _00012_;
  assign mux_303_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_301 : or_528_nl;
  assign mux_301_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_365_cse : or_tmp_522;
  assign mux_300_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_674_nl : nor_675_nl;
  assign mux_299_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_676_nl : nor_677_nl;
  assign mux_297_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_380 : or_tmp_505;
  assign mux_296_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_292 : mux_295_nl;
  assign mux_295_nl = lut_lookup_else_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_505 : mux_294_nl;
  assign mux_294_nl = cfg_lut_le_function_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00010_ : or_tmp_505;
  assign mux_291_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_678_nl : mux_290_nl;
  assign mux_290_nl = lut_lookup_else_if_lor_6_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_679_nl : nor_680_nl;
  assign mux_289_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_681_nl : mux_288_nl;
  assign mux_288_nl = lut_lookup_else_if_lor_6_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_682_nl : nor_683_nl;
  assign mux_287_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_684_nl : nor_685_nl;
  assign mux_286_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_686_nl : nor_687_nl;
  assign mux_1152_nl = cfg_lut_hybrid_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1151_nl : and_451_nl;
  assign mux_1151_nl = cfg_lut_uflow_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1523 : _00011_;
  assign mux_281_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_279 : or_475_nl;
  assign mux_279_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_690_cse : nor_689_nl;
  assign mux_278_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_690_cse : nor_691_nl;
  assign mux_277_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_692_nl : nor_693_nl;
  assign mux_276_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_852_cse : and_843_cse;
  assign mux_274_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_270 : mux_273_nl;
  assign mux_273_nl = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_456 : mux_272_nl;
  assign mux_272_nl = cfg_lut_le_function_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00010_ : or_tmp_456;
  assign mux_270_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_694_nl : nor_695_nl;
  assign mux_269_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_445_nl : or_tmp_447;
  assign mux_268_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_696_nl : nor_697_nl;
  assign mux_267_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_698_nl : nor_699_nl;
  assign mux_1139_nl = cfg_lut_hybrid_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1138_nl : and_447_nl;
  assign mux_1138_nl = cfg_lut_uflow_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1513 : _00009_;
  assign lut_lookup_if_else_else_else_else_mux_3_nl = IsNaN_8U_23U_6_land_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13544|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13543" *) lut_lookup_4_if_else_else_else_else_if_lshift_itm : lut_lookup_4_if_else_else_else_else_else_rshift_itm;
  assign lut_lookup_if_else_else_else_else_mux_2_nl = IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13544|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13543" *) lut_lookup_3_if_else_else_else_else_if_lshift_itm : lut_lookup_3_if_else_else_else_else_else_rshift_itm;
  assign lut_lookup_if_else_else_else_else_mux_1_nl = IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13544|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13543" *) lut_lookup_2_if_else_else_else_else_if_lshift_itm : lut_lookup_2_if_else_else_else_else_else_rshift_itm;
  assign lut_lookup_if_else_else_else_else_mux_nl = IsNaN_8U_23U_6_land_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13544|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13543" *) lut_lookup_1_if_else_else_else_else_if_lshift_itm : lut_lookup_1_if_else_else_else_else_else_rshift_itm;
  assign mux_265_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_80_nl : and_81_nl;
  assign mux_262_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_260_nl : mux_261_nl;
  assign mux_261_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_79_nl : nor_700_nl;
  assign mux_260_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_19 : nor_879_nl;
  assign mux_257_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_705_nl : nor_706_nl;
  assign mux_256_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_254_nl : mux_255_nl;
  assign mux_255_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_312_cse : or_411_nl;
  assign mux_254_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : or_406_nl;
  assign mux_253_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_75_nl : and_76_nl;
  assign mux_250_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_248_nl : mux_249_nl;
  assign mux_249_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_74_nl : _00008_;
  assign mux_248_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_14 : nor_880_nl;
  assign mux_245_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_711_nl : nor_712_nl;
  assign mux_244_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_241_nl : mux_243_nl;
  assign mux_243_nl = lut_lookup_else_else_else_asn_mdf_3_sva_st_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_242_nl : or_tmp_380;
  assign mux_242_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_312_cse : or_tmp_378;
  assign mux_241_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : or_374_nl;
  assign mux_240_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_70_nl : and_71_nl;
  assign mux_237_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_235_nl : mux_236_nl;
  assign mux_236_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_69_nl : nor_714_nl;
  assign mux_235_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_27 : nor_713_nl;
  assign mux_232_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_719_nl : nor_720_nl;
  assign mux_231_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_229_nl : mux_230_nl;
  assign mux_230_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_312_cse : or_346_nl;
  assign mux_229_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : or_341_nl;
  assign mux_228_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_63_nl : and_64_nl;
  assign mux_225_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_223_nl : mux_224_nl;
  assign mux_224_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_62_nl : nor_721_nl;
  assign mux_223_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_5 : nor_881_nl;
  assign mux_219_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_726_nl : nor_727_nl;
  assign mux_218_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_216_nl : mux_217_nl;
  assign mux_217_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_312_cse : or_315_nl;
  assign mux_216_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : or_311_nl;
  assign mux_215_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_213_nl : mux_214_nl;
  assign mux_214_nl = FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : _00004_;
  assign mux_213_nl = IsNaN_8U_23U_7_land_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : _00003_;
  assign mux_211_nl = _03413_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_210_nl : mux_209_nl;
  assign mux_210_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_306_nl : mux_tmp_207;
  assign mux_209_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nand_76_nl : mux_tmp_207;
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_6_nl = FpNormalize_8U_49U_2_oelse_not_15 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl : 8'b00000000;
  assign mux_207_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_204_nl : and_59_nl;
  assign mux_206_nl = cfg_precision_1_sva_st_70[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_57 : mux_205_nl;
  assign mux_205_nl = cfg_precision_1_sva_st_70[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_730_nl : nor_tmp_57;
  assign mux_204_nl = reg_cfg_precision_1_sva_st_13_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_55 : mux_203_nl;
  assign mux_203_nl = reg_cfg_precision_1_sva_st_13_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_729_nl : nor_tmp_55;
  assign mux_202_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_732_nl : nor_733_nl;
  assign mux_200_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_198_nl : mux_199_nl;
  assign mux_199_nl = and_859_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : _00004_;
  assign mux_198_nl = and_858_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : _00003_;
  assign mux_1244_nl = lut_lookup_4_if_else_else_acc_nl[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1995_nl : mux_1243_nl;
  assign mux_1243_nl = reg_cfg_precision_1_sva_st_13_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1707 : mux_1242_nl;
  assign mux_1242_nl = reg_cfg_precision_1_sva_st_13_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00007_ : or_tmp_1707;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_8_nl = FpNormalize_8U_49U_oelse_not_15 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt[5:0] : 6'b000000;
  assign mux_1240_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_4_land_lpi_1_dfm_4 : reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_6_nl = FpNormalize_8U_49U_oelse_not_15 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13510|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13509" *) lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt[7:6] : 2'b00;
  assign mux_1239_nl = _02717_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1238_nl : or_2078_nl;
  assign mux_1238_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1697 : or_1983_nl;
  assign mux_174_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_32_nl : mux_173_nl;
  assign mux_173_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : mux_1212_nl;
  assign mux_1212_nl = FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00001_ : or_tmp_63;
  assign mux_32_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : mux_31_nl;
  assign mux_31_nl = IsNaN_8U_23U_1_land_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00000_ : or_1689_cse;
  assign mux_171_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_169_nl : mux_170_nl;
  assign mux_170_nl = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : _00004_;
  assign mux_169_nl = IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : _00003_;
  assign mux_167_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_165_nl : mux_166_nl;
  assign mux_166_nl = lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : or_251_nl;
  assign mux_165_nl = lut_lookup_3_FpMantRNE_49U_24U_2_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : or_247_nl;
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_4_nl = FpNormalize_8U_49U_2_oelse_not_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl : 8'b00000000;
  assign mux_164_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_161_nl : and_54_nl;
  assign mux_163_nl = cfg_precision_1_sva_st_70[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_46 : mux_162_nl;
  assign mux_162_nl = cfg_precision_1_sva_st_70[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_743_nl : nor_tmp_46;
  assign mux_161_nl = reg_cfg_precision_1_sva_st_13_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_44 : mux_160_nl;
  assign mux_160_nl = reg_cfg_precision_1_sva_st_13_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_742_nl : nor_tmp_44;
  assign mux_159_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_745_nl : nor_746_nl;
  assign mux_157_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_155_nl : mux_156_nl;
  assign mux_156_nl = and_862_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : _00004_;
  assign mux_155_nl = and_861_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : _00003_;
  assign mux_1237_nl = lut_lookup_3_if_else_else_acc_nl[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1976_nl : mux_1236_nl;
  assign mux_1236_nl = reg_cfg_precision_1_sva_st_13_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_48_cse : mux_1235_nl;
  assign mux_1235_nl = reg_cfg_precision_1_sva_st_13_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00006_ : or_48_cse;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_9_nl = FpNormalize_8U_49U_oelse_not_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt[5:0] : 6'b000000;
  assign mux_1233_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_4_land_3_lpi_1_dfm_5 : IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_4_nl = FpNormalize_8U_49U_oelse_not_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13510|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13509" *) lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt[7:6] : 2'b00;
  assign mux_1232_nl = _02693_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1231_nl : or_2079_nl;
  assign mux_1231_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1684 : or_1964_nl;
  assign mux_138_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_27_nl : mux_137_nl;
  assign mux_137_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : mux_1211_nl;
  assign mux_1211_nl = FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00001_ : or_tmp_63;
  assign mux_27_nl = or_48_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : _00000_;
  assign mux_135_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_133_nl : mux_134_nl;
  assign mux_134_nl = FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : _00004_;
  assign mux_133_nl = IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : _00005_;
  assign mux_131_nl = or_tmp_63 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nand_tmp_4 : mux_130_nl;
  assign mux_130_nl = or_184_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_49_nl : nand_tmp_4;
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_2_nl = FpNormalize_8U_49U_2_oelse_not_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl : 8'b00000000;
  assign mux_128_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_125_nl : and_48_nl;
  assign mux_127_nl = cfg_precision_1_sva_st_70[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_34 : mux_126_nl;
  assign mux_126_nl = cfg_precision_1_sva_st_70[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_758_nl : nor_tmp_34;
  assign mux_125_nl = reg_cfg_precision_1_sva_st_13_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_32 : mux_124_nl;
  assign mux_124_nl = reg_cfg_precision_1_sva_st_13_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_757_nl : nor_tmp_32;
  assign mux_123_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_760_nl : nor_761_nl;
  assign mux_121_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_119_nl : mux_120_nl;
  assign mux_120_nl = and_865_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : _00004_;
  assign mux_119_nl = and_864_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : _00003_;
  assign mux_1230_nl = reg_cfg_precision_1_sva_st_13_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1678 : mux_1229_nl;
  assign mux_1229_nl = reg_cfg_precision_1_sva_st_13_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_852_nl : or_tmp_1678;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_10_nl = FpNormalize_8U_49U_oelse_not_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt[5:0] : 6'b000000;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_2_nl = FpNormalize_8U_49U_oelse_not_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13510|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13509" *) lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt[7:6] : 2'b00;
  assign mux_1226_nl = _02672_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1225_nl : or_2080_nl;
  assign mux_1225_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1674 : or_1948_nl;
  assign mux_89_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_23_nl : mux_88_nl;
  assign mux_88_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : mux_87_nl;
  assign mux_87_nl = FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00001_ : or_tmp_63;
  assign mux_23_nl = or_40_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : _00000_;
  assign mux_86_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_84_nl : mux_85_nl;
  assign mux_85_nl = FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : _00004_;
  assign mux_84_nl = IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : _00003_;
  assign mux_82_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_75_nl : mux_81_nl;
  assign mux_81_nl = or_125_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_78 : mux_80_nl;
  assign mux_80_nl = IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00001_ : mux_tmp_78;
  assign mux_75_nl = or_120_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_72 : mux_74_nl;
  assign mux_74_nl = IsNaN_8U_23U_8_land_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00000_ : mux_tmp_72;
  assign mux_69_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_67_nl : mux_68_nl;
  assign mux_68_nl = lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : or_118_nl;
  assign mux_67_nl = lut_lookup_1_FpMantRNE_49U_24U_2_else_and_tmp ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : or_114_nl;
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_nl = FpNormalize_8U_49U_2_oelse_not_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl : 8'b00000000;
  assign mux_66_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_63_nl : and_45_nl;
  assign mux_65_nl = cfg_precision_1_sva_st_70[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_14 : mux_64_nl;
  assign mux_64_nl = cfg_precision_1_sva_st_70[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_770_nl : nor_tmp_14;
  assign mux_63_nl = reg_cfg_precision_1_sva_st_13_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_12 : mux_62_nl;
  assign mux_62_nl = reg_cfg_precision_1_sva_st_13_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_769_nl : nor_tmp_12;
  assign mux_61_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_772_nl : nor_773_nl;
  assign mux_59_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_57_nl : mux_58_nl;
  assign mux_58_nl = and_869_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : _00004_;
  assign mux_57_nl = and_868_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : _00003_;
  assign mux_1224_nl = lut_lookup_1_if_else_else_acc_nl[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1941_nl : mux_1223_nl;
  assign mux_1223_nl = reg_cfg_precision_1_sva_st_13_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1671 : mux_1222_nl;
  assign mux_1222_nl = reg_cfg_precision_1_sva_st_13_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00002_ : or_tmp_1671;
  assign mux_1125_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_dcpl_51 : and_896_cse;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_11_nl = FpNormalize_8U_49U_oelse_not_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt[5:0] : 6'b000000;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_nl = FpNormalize_8U_49U_oelse_not_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13510|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13509" *) lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt[7:6] : 2'b00;
  assign mux_1219_nl = _02652_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1218_nl : or_2081_nl;
  assign mux_1218_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1663 : or_1931_nl;
  assign mux_39_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_13_nl : mux_38_nl;
  assign mux_38_nl = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : mux_1210_nl;
  assign mux_1210_nl = FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00001_ : or_tmp_63;
  assign mux_13_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : mux_1209_nl;
  assign mux_1209_nl = IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00000_ : or_1689_cse;
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_11_nl = FpAdd_8U_23U_b_right_shift_qif_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) _00043_ : _00045_;
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_10_nl = FpAdd_8U_23U_b_right_shift_qif_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) chn_lut_in_rsci_d_mxwt[126:119] : cfg_lut_le_start_rsci_d[30:23];
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_15_nl = FpAdd_8U_23U_b_right_shift_qif_and_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) _00043_ : _00044_;
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_14_nl = FpAdd_8U_23U_b_right_shift_qif_and_tmp_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) chn_lut_in_rsci_d_mxwt[94:87] : cfg_lut_le_start_rsci_d[30:23];
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_13_nl = FpAdd_8U_23U_b_right_shift_qif_and_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) _00043_ : _00042_;
  assign FpAdd_8U_23U_a_right_shift_qelse_mux_12_nl = FpAdd_8U_23U_b_right_shift_qif_and_tmp_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) chn_lut_in_rsci_d_mxwt[62:55] : cfg_lut_le_start_rsci_d[30:23];
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_11_nl = FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) _00041_ : _00040_;
  assign FpAdd_8U_23U_2_a_right_shift_qelse_mux_10_nl = FpAdd_8U_23U_2_b_right_shift_qif_and_tmp_1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) chn_lut_in_rsci_d_mxwt[30:23] : cfg_lut_lo_start_rsci_d[30:23];
  assign lut_lookup_else_2_mux_118_nl = lut_lookup_4_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_lut_lookup_else_2_if_and_6_nl : lut_lookup_else_2_else_mux_76_nl;
  assign lut_lookup_else_2_else_mux_76_nl = _03728_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_56_nl : lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_6_cse;
  assign lut_lookup_else_2_else_else_mux_56_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_6_cse : lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_14_nl;
  assign lut_lookup_else_2_mux_117_nl = lut_lookup_4_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_lut_lookup_else_2_if_and_7_nl : lut_lookup_else_2_else_mux_77_nl;
  assign lut_lookup_else_2_else_mux_77_nl = _03728_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_57_nl : lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_7_cse;
  assign lut_lookup_else_2_else_else_mux_57_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_7_cse : lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_15_nl;
  assign lut_lookup_if_2_mux_24_nl = cfg_lut_uflow_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_mux_116_nl = lut_lookup_4_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) z_out_3 : lut_lookup_else_2_else_mux_78_nl;
  assign lut_lookup_else_2_else_mux_78_nl = _03728_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_58_nl : lut_lookup_else_2_else_if_mux_17_cse_mx0;
  assign lut_lookup_else_2_else_else_mux_58_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_mux_17_cse_mx0 : z_out_3;
  assign lut_lookup_else_2_mux_106_nl = lut_lookup_4_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) cfg_lut_oflow_priority_1_sva_10 : lut_lookup_else_2_else_mux_63_nl;
  assign lut_lookup_else_2_else_mux_63_nl = _03728_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_48_nl : cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_mux_48_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) cfg_lut_hybrid_priority_1_sva_10 : lut_lookup_le_miss_sva;
  assign lut_lookup_else_2_mux_115_nl = lut_lookup_3_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_lut_lookup_else_2_if_and_4_nl : lut_lookup_else_2_else_mux_56_nl;
  assign lut_lookup_else_2_else_mux_56_nl = _03727_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_41_nl : lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_4_cse;
  assign lut_lookup_else_2_else_else_mux_41_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_4_cse : lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_10_nl;
  assign lut_lookup_else_2_mux_114_nl = lut_lookup_3_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_lut_lookup_else_2_if_and_5_nl : lut_lookup_else_2_else_mux_57_nl;
  assign lut_lookup_else_2_else_mux_57_nl = _03727_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_42_nl : lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_5_cse;
  assign lut_lookup_else_2_else_else_mux_42_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_5_cse : lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_11_nl;
  assign lut_lookup_if_2_mux_23_nl = cfg_lut_uflow_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_mux_113_nl = lut_lookup_3_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) z_out_2 : lut_lookup_else_2_else_mux_58_nl;
  assign lut_lookup_else_2_else_mux_58_nl = _03727_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_43_nl : lut_lookup_else_2_else_if_mux_12_cse_mx0;
  assign lut_lookup_else_2_else_else_mux_43_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_mux_12_cse_mx0 : z_out_2;
  assign lut_lookup_else_2_mux_105_nl = lut_lookup_3_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) cfg_lut_oflow_priority_1_sva_10 : lut_lookup_else_2_else_mux_43_nl;
  assign lut_lookup_else_2_else_mux_43_nl = _03727_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_33_nl : cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_mux_33_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_9_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) cfg_lut_hybrid_priority_1_sva_10 : lut_lookup_le_miss_3_sva;
  assign lut_lookup_else_2_mux_112_nl = lut_lookup_2_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_lut_lookup_else_2_if_and_2_nl : lut_lookup_else_2_else_mux_36_nl;
  assign lut_lookup_else_2_else_mux_36_nl = _03726_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_26_nl : lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_2_cse;
  assign lut_lookup_else_2_else_else_mux_26_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_2_cse : lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_6_nl;
  assign lut_lookup_else_2_mux_111_nl = lut_lookup_2_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_lut_lookup_else_2_if_and_3_nl : lut_lookup_else_2_else_mux_37_nl;
  assign lut_lookup_else_2_else_mux_37_nl = _03726_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_27_nl : lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_3_cse;
  assign lut_lookup_else_2_else_else_mux_27_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_3_cse : lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_7_nl;
  assign lut_lookup_if_2_mux_22_nl = cfg_lut_uflow_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_mux_110_nl = lut_lookup_2_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) z_out_1 : lut_lookup_else_2_else_mux_38_nl;
  assign lut_lookup_else_2_else_mux_38_nl = _03726_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_28_nl : lut_lookup_else_2_else_if_mux_7_cse_mx0;
  assign lut_lookup_else_2_else_else_mux_28_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_mux_7_cse_mx0 : z_out_1;
  assign lut_lookup_else_2_mux_104_nl = lut_lookup_2_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) cfg_lut_oflow_priority_1_sva_10 : lut_lookup_else_2_else_mux_23_nl;
  assign lut_lookup_else_2_else_mux_23_nl = _03726_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_18_nl : cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_mux_18_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_5_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) cfg_lut_hybrid_priority_1_sva_10 : lut_lookup_le_miss_2_sva;
  assign lut_lookup_else_2_mux_109_nl = lut_lookup_1_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_lut_lookup_else_2_if_and_nl : lut_lookup_else_2_else_mux_16_nl;
  assign lut_lookup_else_2_else_mux_16_nl = _03725_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_11_nl : lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_cse;
  assign lut_lookup_else_2_else_else_mux_11_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_cse : lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_2_nl;
  assign lut_lookup_else_2_mux_108_nl = lut_lookup_1_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_lut_lookup_else_2_if_and_1_nl : lut_lookup_else_2_else_mux_17_nl;
  assign lut_lookup_else_2_else_mux_17_nl = _03725_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_12_nl : lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_1_cse;
  assign lut_lookup_else_2_else_else_mux_12_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_lut_lookup_else_2_else_if_and_1_cse : lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_3_nl;
  assign lut_lookup_if_2_mux_21_nl = cfg_lut_uflow_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_mux_107_nl = lut_lookup_1_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) z_out : lut_lookup_else_2_else_mux_18_nl;
  assign lut_lookup_else_2_else_mux_18_nl = _03725_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_13_nl : lut_lookup_else_2_else_if_mux_2_cse_mx0;
  assign lut_lookup_else_2_else_else_mux_13_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_if_mux_2_cse_mx0 : z_out;
  assign lut_lookup_else_2_mux_103_nl = lut_lookup_1_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) cfg_lut_oflow_priority_1_sva_10 : lut_lookup_else_2_else_mux_3_nl;
  assign lut_lookup_else_2_else_mux_3_nl = _03725_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_else_else_mux_3_nl : cfg_lut_hybrid_priority_1_sva_10;
  assign lut_lookup_else_2_else_else_mux_3_nl = lut_lookup_else_2_else_else_else_lut_lookup_else_2_else_else_else_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) cfg_lut_hybrid_priority_1_sva_10 : lut_lookup_le_miss_1_sva;
  assign lut_lookup_else_2_mux_79_nl = lut_lookup_4_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_mux_23_nl : lut_lookup_else_2_else_lut_lookup_else_2_else_and_6_nl;
  assign lut_lookup_else_2_else_else_mux_nl = cfg_lut_hybrid_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0 : lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_if_mux_23_nl = cfg_lut_oflow_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0 : lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_mux_53_nl = lut_lookup_3_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_mux_17_nl : lut_lookup_else_2_else_lut_lookup_else_2_else_and_4_nl;
  assign lut_lookup_else_2_else_else_mux_59_nl = cfg_lut_hybrid_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0 : lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_if_mux_17_nl = cfg_lut_oflow_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0 : lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_mux_27_nl = lut_lookup_2_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_mux_11_nl : lut_lookup_else_2_else_lut_lookup_else_2_else_and_2_nl;
  assign lut_lookup_else_2_else_else_mux_60_nl = cfg_lut_hybrid_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0 : lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_if_mux_11_nl = cfg_lut_oflow_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0 : lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_mux_1_nl = lut_lookup_1_else_2_and_svs ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_if_mux_5_nl : lut_lookup_else_2_else_lut_lookup_else_2_else_and_nl;
  assign lut_lookup_else_2_else_else_mux_61_nl = cfg_lut_hybrid_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0 : lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0;
  assign lut_lookup_else_2_if_mux_5_nl = cfg_lut_oflow_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0 : lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0;
  assign mux_tmp_1257 = lut_lookup_else_1_lut_lookup_else_1_and_10_itm_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1261_nl : nor_814_nl;
  assign mux_1261_nl = or_2055_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_unequal_tmp_13 : or_2056_nl;
  assign mux_tmp_1253 = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_1_lut_lookup_else_1_and_7_itm_2 : nor_817_nl;
  assign mux_tmp_1250 = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_1_lut_lookup_else_1_and_4_itm_2 : nor_820_nl;
  assign mux_tmp_1247 = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_1_lut_lookup_else_1_and_1_itm_2 : nor_823_nl;
  assign mux_1241_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1991_nl : or_1992_nl;
  assign mux_1234_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1972_nl : or_1973_nl;
  assign mux_1180_nl = cfg_lut_hybrid_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_438_nl : mux_1179_nl;
  assign mux_1179_nl = cfg_lut_uflow_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00013_ : or_tmp_1545;
  assign mux_1167_nl = cfg_lut_hybrid_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_440_nl : mux_1166_nl;
  assign mux_1166_nl = cfg_lut_uflow_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00012_ : or_tmp_1534;
  assign mux_1154_nl = cfg_lut_hybrid_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_442_nl : mux_1153_nl;
  assign mux_1153_nl = cfg_lut_uflow_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00011_ : or_tmp_1523;
  assign mux_1141_nl = cfg_lut_hybrid_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_444_nl : mux_1140_nl;
  assign mux_1140_nl = cfg_lut_uflow_priority_1_sva_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00009_ : or_tmp_1513;
  assign mux_tmp_1175 = lut_lookup_lo_uflow_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_1169 : _00039_;
  assign mux_tmp_1169 = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_129_itm_2 : mux_1168_nl;
  assign mux_1168_nl = or_1202_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_else_lut_lookup_if_else_or_3_cse : or_1618_nl;
  assign mux_tmp_1162 = lut_lookup_lo_uflow_3_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_1156 : _00038_;
  assign mux_tmp_1156 = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_86_itm_2 : mux_1155_nl;
  assign mux_1155_nl = or_1202_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_else_lut_lookup_if_else_or_2_cse : or_1606_nl;
  assign mux_tmp_1149 = lut_lookup_lo_uflow_2_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_1143 : _00037_;
  assign mux_tmp_1143 = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_43_itm_2 : mux_1142_nl;
  assign mux_1142_nl = or_1202_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_else_lut_lookup_if_else_or_1_cse : or_1594_nl;
  assign mux_tmp_1136 = lut_lookup_lo_uflow_1_lpi_1_dfm_3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_1130 : _00036_;
  assign mux_tmp_1130 = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_itm_2 : mux_1129_nl;
  assign mux_1129_nl = or_1202_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_else_lut_lookup_if_else_or_cse : or_1583_nl;
  assign mux_tmp_1101 = or_26_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_1 : not_tmp_422;
  assign mux_tmp_978 = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_826_cse : and_852_cse;
  assign mux_793_cse = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : and_tmp_6;
  assign mux_tmp_704 = cfg_precision_1_sva_st_70[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : nor_622_nl;
  assign mux_tmp_655 = reg_cfg_precision_1_sva_st_13_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : nor_641_nl;
  assign mux_tmp_643 = or_1688_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : mux_639_nl;
  assign mux_639_nl = or_856_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : _00000_;
  assign mux_tmp_618 = or_832_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_617 : nor_647_nl;
  assign mux_tmp_617 = or_841_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00034_ : mux_617_nl;
  assign mux_617_nl = reg_cfg_precision_1_sva_st_13_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00035_ : _00034_;
  assign mux_616_nl = lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_843 : mux_615_nl;
  assign mux_615_nl = FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_874_cse : or_tmp_843;
  assign mux_tmp_596 = or_tmp_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_595 : or_1860_nl;
  assign mux_tmp_595 = _03374_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : _00003_;
  assign mux_595_itm = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_6 : mux_594_nl;
  assign mux_594_nl = reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nand_95_cse : or_1688_cse;
  assign mux_582_itm = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_6 : mux_581_nl;
  assign mux_581_nl = reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nand_95_cse : or_1688_cse;
  assign mux_tmp_475 = _03401_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : _00003_;
  assign mux_tmp_292 = lut_lookup_else_unequal_tmp_12 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_380 : mux_292_nl;
  assign mux_292_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00032_ : or_tmp_380;
  assign mux_tmp_281 = lut_lookup_else_unequal_tmp_18 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_312_cse : _00032_;
  assign mux_tmp_270 = or_1853_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_380 : _00032_;
  assign mux_tmp_265 = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : main_stage_v_5;
  assign mux_tmp_220 = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : main_stage_v_4;
  assign mux_tmp_207 = lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : or_302_nl;
  assign mux_tmp_128 = or_186_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nand_93_nl : or_191_nl;
  assign mux_tmp_78 = or_126_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_76 : mux_78_nl;
  assign mux_78_nl = IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00001_ : mux_tmp_76;
  assign mux_tmp_76 = or_127_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_129 : mux_76_nl;
  assign mux_76_nl = IsNaN_8U_23U_8_land_3_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00001_ : or_tmp_129;
  assign mux_tmp_72 = or_121_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_70 : mux_72_nl;
  assign mux_72_nl = IsNaN_8U_23U_8_land_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00000_ : mux_tmp_70;
  assign mux_tmp_70 = or_122_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_124 : mux_70_nl;
  assign mux_70_nl = IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00000_ : or_tmp_124;
  assign mux_tmp_35 = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : main_stage_v_3;
  assign mux_26_itm = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1688_cse : or_tmp_44;
  assign mux_25_itm = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1688_cse : or_1689_cse;
  assign mux_20_itm = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_8 : or_1689_cse;
  assign not_tmp_47 = or_26_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_779_nl : mux_18_nl;
  assign mux_18_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_1 : _00003_;
  assign mux_tmp_10 = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_1 : main_stage_v_2;
  assign mux_tmp_4 = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_6 : or_1688_cse;
  assign mux_3_itm = or_26_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_4_nl : mux_2_nl;
  assign mux_2_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_6 : _00033_;
  assign lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp = lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[135:127];
  assign FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_2_int_mant_p1_sva_3[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) { 1'b1, FpAdd_8U_23U_2_int_mant_p1_sva_3[48:1] } : FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_7_nl;
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_7_nl = FpNormalize_8U_49U_2_oelse_not_15 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_sva = lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[135:127];
  assign FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_1_int_mant_p1_sva_3[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) { 1'b1, FpAdd_8U_23U_1_int_mant_p1_sva_3[48:1] } : FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl = FpNormalize_8U_49U_oelse_not_15 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) lut_lookup_4_FpNormalize_8U_49U_else_lshift_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp = lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[135:127];
  assign FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_2_int_mant_p1_3_sva_3[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) { 1'b1, FpAdd_8U_23U_2_int_mant_p1_3_sva_3[48:1] } : FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_5_nl;
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_5_nl = FpNormalize_8U_49U_2_oelse_not_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_3_sva = lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[135:127];
  assign FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) { 1'b1, FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:1] } : FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl = FpNormalize_8U_49U_oelse_not_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) lut_lookup_3_FpNormalize_8U_49U_else_lshift_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp = lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[135:127];
  assign FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_2_int_mant_p1_2_sva_3[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) { 1'b1, FpAdd_8U_23U_2_int_mant_p1_2_sva_3[48:1] } : FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_3_nl;
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_3_nl = FpNormalize_8U_49U_2_oelse_not_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_2_sva = lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[135:127];
  assign FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) { 1'b1, FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:1] } : FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl = FpNormalize_8U_49U_oelse_not_11 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) lut_lookup_2_FpNormalize_8U_49U_else_lshift_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp = lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_1_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm[135:127];
  assign FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_2_int_mant_p1_1_sva_3[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) { 1'b1, FpAdd_8U_23U_2_int_mant_p1_1_sva_3[48:1] } : FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_1_nl;
  assign FpNormalize_8U_49U_2_FpNormalize_8U_49U_2_and_1_nl = FpNormalize_8U_49U_2_oelse_not_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign IntSignedShiftRightTZ_32U_8U_9U_ac_int_cctor_1_sva = lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_obits_fixed_or_1_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm[135:127];
  assign FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0 = FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) { 1'b1, FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:1] } : FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl = FpNormalize_8U_49U_oelse_not_9 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) lut_lookup_1_FpNormalize_8U_49U_else_lshift_itm : 49'b0000000000000000000000000000000000000000000000000;
  assign FpAdd_8U_23U_2_a_right_shift_qr_lpi_1_dfm = FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) 8'b00000000 : FpAdd_8U_23U_2_a_right_shift_qr_sva_3;
  assign FpAdd_8U_23U_2_b_right_shift_qr_lpi_1_dfm = FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) FpAdd_8U_23U_2_a_right_shift_qr_sva_3 : 8'b00000000;
  assign FpAdd_8U_23U_2_addend_smaller_qr_lpi_1_dfm_mx0 = FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_2_addend_larger_asn_1_mx0w1 : FpAdd_8U_23U_2_a_int_mant_p1_sva;
  assign FpAdd_8U_23U_2_addend_larger_qr_lpi_1_dfm_mx0 = FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_2_a_int_mant_p1_sva : FpAdd_8U_23U_2_addend_larger_asn_1_mx0w1;
  assign FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1 : FpAdd_8U_23U_1_a_int_mant_p1_sva;
  assign FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_1_a_int_mant_p1_sva : FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1;
  assign FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm = FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) 8'b00000000 : FpAdd_8U_23U_1_a_right_shift_qr_sva_3;
  assign FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm = FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) FpAdd_8U_23U_1_a_right_shift_qr_sva_3 : 8'b00000000;
  assign FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_addend_larger_asn_1_mx0w1 : FpAdd_8U_23U_a_int_mant_p1_sva;
  assign FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_a_int_mant_p1_sva : FpAdd_8U_23U_addend_larger_asn_1_mx0w1;
  assign FpAdd_8U_23U_2_a_right_shift_qr_3_lpi_1_dfm = FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) 8'b00000000 : FpAdd_8U_23U_2_a_right_shift_qr_3_sva_3;
  assign FpAdd_8U_23U_2_b_right_shift_qr_3_lpi_1_dfm = FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) FpAdd_8U_23U_2_a_right_shift_qr_3_sva_3 : 8'b00000000;
  assign FpAdd_8U_23U_2_addend_smaller_qr_3_lpi_1_dfm_mx0 = FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_2_addend_larger_asn_7_mx0w1 : FpAdd_8U_23U_2_a_int_mant_p1_3_sva;
  assign FpAdd_8U_23U_2_addend_larger_qr_3_lpi_1_dfm_mx0 = FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_2_a_int_mant_p1_3_sva : FpAdd_8U_23U_2_addend_larger_asn_7_mx0w1;
  assign FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1 : FpAdd_8U_23U_1_a_int_mant_p1_3_sva;
  assign FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_1_a_int_mant_p1_3_sva : FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1;
  assign FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm = FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) 8'b00000000 : FpAdd_8U_23U_1_a_right_shift_qr_3_sva_3;
  assign FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm = FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) FpAdd_8U_23U_1_a_right_shift_qr_3_sva_3 : 8'b00000000;
  assign FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_addend_larger_asn_7_mx0w1 : FpAdd_8U_23U_a_int_mant_p1_3_sva;
  assign FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_a_int_mant_p1_3_sva : FpAdd_8U_23U_addend_larger_asn_7_mx0w1;
  assign FpAdd_8U_23U_2_a_right_shift_qr_2_lpi_1_dfm = FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) 8'b00000000 : FpAdd_8U_23U_2_a_right_shift_qr_2_sva_3;
  assign FpAdd_8U_23U_2_b_right_shift_qr_2_lpi_1_dfm = FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) FpAdd_8U_23U_2_a_right_shift_qr_2_sva_3 : 8'b00000000;
  assign FpAdd_8U_23U_2_addend_smaller_qr_2_lpi_1_dfm_mx0 = FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_2_addend_larger_asn_13_mx0w1 : FpAdd_8U_23U_2_a_int_mant_p1_2_sva;
  assign FpAdd_8U_23U_2_addend_larger_qr_2_lpi_1_dfm_mx0 = FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_2_a_int_mant_p1_2_sva : FpAdd_8U_23U_2_addend_larger_asn_13_mx0w1;
  assign FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1 : FpAdd_8U_23U_1_a_int_mant_p1_2_sva;
  assign FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_1_a_int_mant_p1_2_sva : FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1;
  assign FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm = FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) 8'b00000000 : FpAdd_8U_23U_1_a_right_shift_qr_2_sva_3;
  assign FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm = FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) FpAdd_8U_23U_1_a_right_shift_qr_2_sva_3 : 8'b00000000;
  assign FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_addend_larger_asn_13_mx0w1 : FpAdd_8U_23U_a_int_mant_p1_2_sva;
  assign FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_a_int_mant_p1_2_sva : FpAdd_8U_23U_addend_larger_asn_13_mx0w1;
  assign FpAdd_8U_23U_2_a_right_shift_qr_1_lpi_1_dfm = FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) 8'b00000000 : FpAdd_8U_23U_2_a_right_shift_qr_1_sva_3;
  assign FpAdd_8U_23U_2_b_right_shift_qr_1_lpi_1_dfm = FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) FpAdd_8U_23U_2_a_right_shift_qr_1_sva_3 : 8'b00000000;
  assign FpAdd_8U_23U_2_addend_smaller_qr_1_lpi_1_dfm_mx0 = FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_2_addend_larger_asn_19_mx0w1 : FpAdd_8U_23U_2_a_int_mant_p1_1_sva;
  assign FpAdd_8U_23U_2_addend_larger_qr_1_lpi_1_dfm_mx0 = FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_2_a_int_mant_p1_1_sva : FpAdd_8U_23U_2_addend_larger_asn_19_mx0w1;
  assign FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1 : FpAdd_8U_23U_1_a_int_mant_p1_1_sva;
  assign FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_1_a_int_mant_p1_1_sva : FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1;
  assign FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm = FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) 8'b00000000 : FpAdd_8U_23U_1_a_right_shift_qr_1_sva_3;
  assign FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm = FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) FpAdd_8U_23U_1_a_right_shift_qr_1_sva_3 : 8'b00000000;
  assign FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_addend_larger_asn_19_mx0w1 : FpAdd_8U_23U_a_int_mant_p1_1_sva;
  assign FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_mx0 = FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13561|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13560" *) FpAdd_8U_23U_a_int_mant_p1_1_sva : FpAdd_8U_23U_addend_larger_asn_19_mx0w1;
  assign _00061_ = IsNaN_8U_23U_10_land_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_3_nl;
  assign _00060_ = lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2[8:0];
  assign _00059_ = IsNaN_8U_23U_6_land_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_3_nl;
  assign _00058_ = lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_sva_2[8:0];
  assign lut_lookup_else_2_else_if_mux_17_cse_mx0 = cfg_lut_hybrid_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0;
  assign lut_lookup_lo_index_0_7_0_lpi_1_dfm_4_mx0_7_6 = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13510|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13509" *) lut_lookup_lo_index_0_7_0_lpi_1_dfm_13[7:6] : lut_lookup_lo_index_0_7_0_lpi_1_dfm_1[7:6];
  assign lut_lookup_le_index_0_6_lpi_1_dfm_8_mx0 = cfg_lut_le_function_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_178_nl : lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2;
  assign lut_lookup_else_mux_178_nl = lut_lookup_else_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2 : lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_3_nl;
  assign lut_lookup_lo_index_0_8_lpi_1_dfm_2_mx0 = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_1_lut_lookup_else_1_and_10_itm_2 : lut_lookup_if_1_lut_lookup_if_1_and_14_nl;
  assign _00057_ = IsNaN_8U_23U_10_land_3_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_2_nl;
  assign _00056_ = lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2[8:0];
  assign _00055_ = IsNaN_8U_23U_6_land_3_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_2_nl;
  assign _00054_ = lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_3_sva_2[8:0];
  assign lut_lookup_else_2_else_if_mux_12_cse_mx0 = cfg_lut_hybrid_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0;
  assign lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_4_mx0_7_6 = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13510|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13509" *) lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_13[7:6] : lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_1[7:6];
  assign lut_lookup_lo_index_0_8_3_lpi_1_dfm_2_mx0 = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_1_lut_lookup_else_1_and_7_itm_2 : lut_lookup_if_1_lut_lookup_if_1_and_13_nl;
  assign lut_lookup_le_index_0_6_3_lpi_1_dfm_8_mx0 = cfg_lut_le_function_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_176_nl : lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2;
  assign lut_lookup_else_mux_176_nl = lut_lookup_else_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2 : lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_2_nl;
  assign _00053_ = IsNaN_8U_23U_10_land_2_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_1_nl;
  assign _00052_ = lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2[8:0];
  assign _00051_ = IsNaN_8U_23U_6_land_2_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_1_nl;
  assign _00050_ = lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_2_sva_2[8:0];
  assign lut_lookup_else_2_else_if_mux_7_cse_mx0 = cfg_lut_hybrid_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0;
  assign lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_4_mx0_7_6 = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13510|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13509" *) lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_13[7:6] : lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_1[7:6];
  assign lut_lookup_lo_index_0_8_2_lpi_1_dfm_2_mx0 = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_1_lut_lookup_else_1_and_4_itm_2 : lut_lookup_if_1_lut_lookup_if_1_and_12_nl;
  assign lut_lookup_le_index_0_6_2_lpi_1_dfm_8_mx0 = cfg_lut_le_function_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_174_nl : lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2;
  assign lut_lookup_else_mux_174_nl = lut_lookup_else_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2 : lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_1_nl;
  assign _00049_ = IsNaN_8U_23U_10_land_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_nor_nl;
  assign _00048_ = lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2[8:0];
  assign _00047_ = IsNaN_8U_23U_6_land_1_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_nor_nl;
  assign _00046_ = lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) 9'b111111111 : FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_1_sva_2[8:0];
  assign lut_lookup_else_2_else_if_mux_2_cse_mx0 = cfg_lut_hybrid_priority_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6[0] : lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0;
  assign lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_4_mx0_7_6 = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13510|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13509" *) lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_13[7:6] : lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_1[7:6];
  assign lut_lookup_lo_index_0_8_1_lpi_1_dfm_2_mx0 = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_1_lut_lookup_else_1_and_1_itm_2 : lut_lookup_if_1_lut_lookup_if_1_and_11_nl;
  assign lut_lookup_le_index_0_6_1_lpi_1_dfm_8_mx0 = cfg_lut_le_function_1_sva_10 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_172_nl : lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2;
  assign lut_lookup_else_mux_172_nl = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2 : lut_lookup_else_if_lut_lookup_else_if_lut_lookup_else_if_nor_nl;
  assign FpAdd_8U_23U_2_o_mant_lpi_1_dfm_2_mx0 = IsNaN_8U_23U_7_land_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) lut_in_data_sva_156[118:96] : FpAdd_8U_23U_2_asn_35_mx0w1;
  assign FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0 = lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_7_nl : FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5;
  assign FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx0 = IsNaN_8U_23U_3_land_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) lut_in_data_sva_156[118:96] : FpAdd_8U_23U_asn_35_mx0w1;
  assign FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0 = reg_lut_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_7_nl : FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6;
  assign FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_2_mx0 = IsNaN_8U_23U_7_land_3_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) lut_in_data_sva_156[86:64] : FpAdd_8U_23U_2_asn_40_mx0w1;
  assign FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0 = lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_6_nl : FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5;
  assign FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx0 = IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) lut_in_data_sva_156[86:64] : FpAdd_8U_23U_asn_40_mx0w1;
  assign FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0 = reg_lut_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_6_nl : FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6;
  assign FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_2_mx0 = IsNaN_8U_23U_7_land_2_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) lut_in_data_sva_156[54:32] : FpAdd_8U_23U_2_asn_45_mx0w1;
  assign FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0 = lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_5_nl : FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5;
  assign FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx0 = IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) lut_in_data_sva_156[54:32] : FpAdd_8U_23U_asn_45_mx0w1;
  assign FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0 = reg_lut_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_5_nl : FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6;
  assign FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_2_mx0 = IsNaN_8U_23U_7_land_1_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) lut_in_data_sva_156[22:0] : FpAdd_8U_23U_2_asn_50_mx0w1;
  assign FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0 = lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_if_4_FpAdd_8U_23U_2_if_4_or_4_nl : FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5;
  assign FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx0 = IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) lut_in_data_sva_156[22:0] : FpAdd_8U_23U_asn_50_mx0w1;
  assign FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0 = reg_lut_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_4_nl : FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6;
  assign FpAdd_8U_23U_2_asn_35_mx0w1 = IsNaN_8U_23U_8_land_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) cfg_lut_lo_start_1_sva_3_30_0_1[22:0] : FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_7_nl;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_7_nl = FpAdd_8U_23U_2_is_inf_lpi_1_dfm_2_mx0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) 23'b11111111111111111111111 : lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl;
  assign FpAdd_8U_23U_asn_35_mx0w1 = IsNaN_8U_23U_1_land_lpi_1_dfm_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) cfg_lut_le_start_1_sva_3_30_0_1[22:0] : FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl;
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_7_nl = FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) 23'b11111111111111111111111 : lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl;
  assign FpAdd_8U_23U_2_asn_40_mx0w1 = IsNaN_8U_23U_8_land_3_lpi_1_dfm_5 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) cfg_lut_lo_start_1_sva_3_30_0_1[22:0] : FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_6_nl;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_6_nl = FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_2_mx0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) 23'b11111111111111111111111 : lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl;
  assign FpAdd_8U_23U_asn_40_mx0w1 = IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) cfg_lut_le_start_1_sva_3_30_0_1[22:0] : FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl;
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_6_nl = FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) 23'b11111111111111111111111 : lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl;
  assign FpAdd_8U_23U_2_asn_45_mx0w1 = IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) cfg_lut_lo_start_1_sva_3_30_0_1[22:0] : FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_5_nl;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_5_nl = FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_2_mx0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) 23'b11111111111111111111111 : lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl;
  assign FpAdd_8U_23U_asn_45_mx0w1 = IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) cfg_lut_le_start_1_sva_3_30_0_1[22:0] : FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl;
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_5_nl = FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) 23'b11111111111111111111111 : lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl;
  assign FpAdd_8U_23U_2_asn_50_mx0w1 = IsNaN_8U_23U_8_land_2_lpi_1_dfm_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) cfg_lut_lo_start_1_sva_3_30_0_1[22:0] : FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_4_nl;
  assign FpAdd_8U_23U_2_FpAdd_8U_23U_2_or_4_nl = FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_2_mx0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) 23'b11111111111111111111111 : lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl;
  assign FpAdd_8U_23U_asn_50_mx0w1 = IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) cfg_lut_le_start_1_sva_3_30_0_1[22:0] : FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl;
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_4_nl = FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) 23'b11111111111111111111111 : lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl;
  assign lut_lookup_if_mux_mx0w1 = _02050_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_if_lut_lookup_if_if_or_nl : lut_lookup_if_else_lut_lookup_if_else_or_cse;
  assign lut_lookup_if_mux_41_mx0w1 = _02050_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_if_lut_lookup_if_if_or_1_nl : lut_lookup_if_else_lut_lookup_if_else_or_1_cse;
  assign lut_lookup_if_mux_82_mx0w1 = _02050_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_if_lut_lookup_if_if_or_2_nl : lut_lookup_if_else_lut_lookup_if_else_or_2_cse;
  assign lut_lookup_if_mux_123_mx0w1 = _02050_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_if_lut_lookup_if_if_or_3_nl : lut_lookup_if_else_lut_lookup_if_else_or_3_cse;
  assign mux_1115_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_178 : mux_tmp_1104;
  assign mux_1106_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_1104 : and_42_cse;
  assign mux_1074_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_465_nl : nor_466_nl;
  assign mux_1067_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_478_nl : nor_479_nl;
  assign mux_1056_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_42_cse : mux_tmp_704;
  assign mux_1053_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_42_cse : and_tmp_6;
  assign mux_1004_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_178_cse : and_1179_nl;
  assign mux_982_cse = or_66_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_2 : and_42_cse;
  assign mux_1269_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : and_164_nl;
  assign mux_1205_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_412_nl : nor_413_nl;
  assign mux_1204_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_414_nl : nor_415_nl;
  assign IntLog2_32U_IntLog2_32U_mux_2_rgt = mux_1187_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13527|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13526" *) lut_lookup_4_IntLog2_32U_and_nl : { 8'b00000000, lut_lookup_lut_lookup_mux_4_nl };
  assign lut_lookup_lut_lookup_mux_4_nl = and_672_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) FpAdd_8U_23U_asn_35_mx0w1 : lut_in_data_sva_156[118:96];
  assign mux_919_nl = lut_lookup_else_unequal_tmp_18 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_917_nl : mux_918_nl;
  assign mux_918_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_6 : and_tmp_83;
  assign mux_917_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) and_tmp_6 : main_stage_v_4;
  assign mux_1278_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : and_153_nl;
  assign mux_1200_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_418_nl : nor_419_nl;
  assign mux_1199_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_420_nl : nor_421_nl;
  assign IntLog2_32U_IntLog2_32U_mux_1_rgt = mux_1187_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13527|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13526" *) lut_lookup_3_IntLog2_32U_and_nl : { 8'b00000000, lut_lookup_lut_lookup_mux_3_nl };
  assign lut_lookup_lut_lookup_mux_3_nl = and_665_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) FpAdd_8U_23U_asn_40_mx0w1 : lut_in_data_sva_156[86:64];
  assign mux_853_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_851_cse : mux_852_nl;
  assign mux_852_nl = and_811_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : and_134_cse;
  assign mux_851_cse = cfg_lut_le_function_1_sva_st_41 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_793_cse : and_826_cse;
  assign mux_1279_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : and_143_nl;
  assign mux_1195_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_424_nl : nor_425_nl;
  assign mux_1194_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_426_nl : nor_427_nl;
  assign IntLog2_32U_IntLog2_32U_mux_rgt = mux_1187_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13527|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13526" *) lut_lookup_2_IntLog2_32U_and_nl : { 8'b00000000, lut_lookup_lut_lookup_mux_nl };
  assign lut_lookup_lut_lookup_mux_nl = and_657_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) FpAdd_8U_23U_asn_45_mx0w1 : lut_in_data_sva_156[54:32];
  assign mux_805_cse = lut_lookup_else_unequal_tmp_18 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : and_tmp_83;
  assign lut_lookup_else_1_else_else_mux1h_1_itm = mux_1187_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13629|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13628" *) lut_lookup_1_else_1_else_else_acc_nl : { 1'b0, FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl };
  assign mux_1280_nl = or_1857_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : and_132_nl;
  assign mux_1190_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_430_nl : nor_431_nl;
  assign mux_1189_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_432_nl : nor_433_nl;
  assign mux_1188_cse = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_434_nl : nor_435_nl;
  assign IntLog2_32U_mux1h_1_itm = mux_1187_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13527|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13526" *) lut_lookup_1_IntLog2_32U_and_nl : { 8'b00000000, lut_lookup_lut_lookup_mux_17_nl };
  assign lut_lookup_lut_lookup_mux_17_nl = and_649_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) FpAdd_8U_23U_asn_50_mx0w1 : lut_in_data_sva_156[22:0];
  assign mux_1187_cse = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1857_cse : or_tmp_314;
  assign mux_775_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_771_cse : mux_774_nl;
  assign mux_774_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_612_cse : mux_773_nl;
  assign mux_773_nl = cfg_precision_1_sva_st_71[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : mux_772_nl;
  assign mux_772_nl = cfg_precision_1_sva_st_71[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_609_nl : main_stage_v_4;
  assign mux_1281_nl = cfg_precision_1_sva_st_70[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_3 : mux_769_nl;
  assign mux_769_nl = cfg_precision_1_sva_st_70[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_606_nl : main_stage_v_3;
  assign mux_755_cse = cfg_precision_1_sva_st_71[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : mux_754_nl;
  assign mux_754_nl = cfg_precision_1_sva_st_71[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00027_ : main_stage_v_4;
  assign mux_749_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_745_cse : mux_748_nl;
  assign mux_748_nl = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_978_cse : mux_747_nl;
  assign mux_747_nl = cfg_precision_1_sva_st_71[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_980 : mux_746_nl;
  assign mux_746_nl = cfg_precision_1_sva_st_71[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00032_ : or_tmp_980;
  assign mux_1282_nl = cfg_precision_1_sva_st_70[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_976 : mux_743_nl;
  assign mux_743_nl = cfg_precision_1_sva_st_70[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00001_ : or_tmp_976;
  assign mux_735_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1285_cse : mux_tmp_281;
  assign mux_729_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_704 : nor_tmp_112;
  assign mux_717_nl = lut_lookup_else_unequal_tmp_18 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_715_nl : mux_716_nl;
  assign mux_716_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1285_cse : _00032_;
  assign mux_715_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_1285_cse : or_312_cse;
  assign mux_707_nl = lut_lookup_else_unequal_tmp_18 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_706_nl : and_120_nl;
  assign mux_706_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_704 : main_stage_v_4;
  assign mux_671_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_670_cse : mux_tmp_292;
  assign mux_1285_cse = cfg_precision_1_sva_st_70[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_63 : mux_668_nl;
  assign mux_668_nl = cfg_precision_1_sva_st_70[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00001_ : or_tmp_63;
  assign mux_1186_nl = reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1696_nl : and_nl;
  assign mux_1185_nl = reg_cfg_lut_le_function_1_sva_st_19_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_6 : IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
  assign mux_580_cse = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) chn_lut_in_rsci_bawt : main_stage_v_1;
  assign mux_366_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_tmp_112 : and_832_cse;
  assign mux_360_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_358_nl : mux_359_nl;
  assign mux_359_nl = lut_lookup_else_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_5 : not_tmp_334;
  assign mux_358_nl = lut_lookup_else_unequal_tmp_12 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : nor_612_cse;
  assign mux_357_nl = lut_lookup_else_unequal_tmp_18 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_356_nl : nor_657_nl;
  assign mux_356_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) main_stage_v_4 : and_832_cse;
  assign lut_lookup_else_mux_186_cse = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_129_itm_2 : lut_lookup_if_mux_123_mx0w1;
  assign mux_330_nl = lut_lookup_else_unequal_tmp_18 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_328_nl : mux_329_nl;
  assign mux_329_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _00032_ : mux_283_cse;
  assign mux_328_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_312_cse : mux_283_cse;
  assign mux_316_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_292 : mux_315_nl;
  assign mux_315_nl = lut_lookup_else_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_456 : mux_272_nl;
  assign lut_lookup_else_mux_184_cse = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_86_itm_2 : lut_lookup_if_mux_82_mx0w1;
  assign lut_lookup_else_mux_182_cse = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_43_itm_2 : lut_lookup_if_mux_41_mx0w1;
  assign mux_285_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_312_cse : or_tmp_478;
  assign mux_284_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) mux_tmp_281 : mux_283_cse;
  assign mux_283_cse = lut_lookup_unequal_tmp_13 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_478 : _00010_;
  assign mux_275_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_380 : or_tmp_456;
  assign lut_lookup_else_mux_180_cse = cfg_lut_le_function_1_sva_st_42 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_itm_2 : lut_lookup_if_mux_mx0w1;
  assign mux_263_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_427 : or_tmp_428;
  assign mux_259_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_701_nl : nor_702_nl;
  assign mux_251_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_395 : or_tmp_397;
  assign mux_247_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_707_nl : nor_708_nl;
  assign mux_238_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_363 : or_365_cse;
  assign mux_234_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_715_nl : nor_716_nl;
  assign mux_226_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_331 : or_332_nl;
  assign mux_222_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_722_nl : nor_723_nl;
  assign mux_220_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_724_nl : nor_725_nl;
  assign mux_177_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_737_nl : nor_738_nl;
  assign mux_141_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_749_nl : nor_750_nl;
  assign mux_132_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_44 : or_tmp_63;
  assign mux_1126_cse = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_dcpl_57 : and_896_cse;
  assign mux_1227_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_4_land_2_lpi_1_dfm_5 : IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5;
  assign mux_92_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_764_nl : nor_765_nl;
  assign mux_83_cse = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_1689_cse : or_tmp_63;
  assign mux_1220_nl = reg_cfg_lut_le_function_1_sva_st_20_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_4_land_1_lpi_1_dfm_4 : IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5;
  assign mux_42_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_775_nl : nor_776_nl;
  assign FpAdd_8U_23U_1_mux1h_7_itm = mux_1122_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) { 2'b00, libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_7 } : FpAdd_8U_23U_1_qr_lpi_1_dfm_5;
  assign FpAdd_8U_23U_1_mux1h_5_itm = mux_1122_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) { 2'b00, libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_6 } : FpAdd_8U_23U_1_qr_4_lpi_1_dfm_5;
  assign FpAdd_8U_23U_1_mux1h_3_itm = mux_1122_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) { 2'b00, libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_5 } : FpAdd_8U_23U_1_qr_3_lpi_1_dfm_5;
  assign mux_1122_cse = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_26_cse : or_66_cse;
  assign FpAdd_8U_23U_1_mux1h_1_itm = mux_1121_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) { 2'b00, libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_4 } : FpAdd_8U_23U_1_qr_2_lpi_1_dfm_5;
  assign mux_1121_nl = reg_cfg_precision_1_sva_st_12_cse_1[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_1490 : mux_1120_nl;
  assign mux_1120_nl = reg_cfg_precision_1_sva_st_12_cse_1[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) nor_783_nl : or_tmp_1490;
  assign mux_4_nl = or_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_tmp_6 : or_tmp_8;
  assign _00471_ = _01136_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11685" *) lut_lookup_1_else_1_acc_nl[32] : lut_lookup_else_1_slc_32_mdf_1_sva_5;
  assign _00475_ = lut_lookup_else_1_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11675" *) lut_lookup_2_else_1_acc_nl[32] : lut_lookup_else_1_slc_32_mdf_2_sva_5;
  assign _00479_ = lut_lookup_else_1_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11675" *) lut_lookup_3_else_1_acc_nl[32] : lut_lookup_else_1_slc_32_mdf_3_sva_5;
  assign _00483_ = lut_lookup_else_1_and_16_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11675" *) lut_lookup_4_else_1_acc_nl[32] : lut_lookup_else_1_slc_32_mdf_sva_5;
  assign _00484_ = _01135_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11665" *) lut_lookup_else_1_slc_32_mdf_sva_5 : lut_lookup_else_1_slc_32_mdf_sva_6;
  assign _00569_ = _01134_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11657" *) lut_lookup_if_else_else_le_data_sub_sva_mx0w0[30:0] : lut_lookup_if_else_else_le_data_sub_sva_1_30_0_1;
  assign _00568_ = _01133_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11649" *) lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0[30:0] : lut_lookup_if_else_else_le_data_sub_3_sva_1_30_0_1;
  assign _00476_ = lut_lookup_else_1_and_13_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11640" *) lut_lookup_else_1_slc_32_mdf_2_sva_5 : lut_lookup_else_1_slc_32_mdf_2_sva_6;
  assign _00480_ = lut_lookup_else_1_and_13_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11640" *) lut_lookup_else_1_slc_32_mdf_3_sva_5 : lut_lookup_else_1_slc_32_mdf_3_sva_6;
  assign _00567_ = _01132_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11631" *) lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0[30:0] : lut_lookup_if_else_else_le_data_sub_2_sva_1_30_0_1;
  assign _00472_ = _01131_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11623" *) lut_lookup_else_1_slc_32_mdf_1_sva_5 : lut_lookup_else_1_slc_32_mdf_1_sva_6;
  assign _00566_ = _01130_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11615" *) lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0[30:0] : lut_lookup_if_else_else_le_data_sub_1_sva_1_30_0_1;
  assign _00466_ = _01129_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11607" *) lut_lookup_else_1_lo_index_u_sva_3 : lut_lookup_else_1_lo_index_u_sva_4;
  assign _00510_ = _01128_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11599" *) lut_lookup_else_else_else_le_index_u_sva_3 : lut_lookup_else_else_else_le_index_u_sva_4;
  assign _00857_ = and_dcpl_148 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_else_else_else_lut_lookup_else_else_else_and_7_nl : lut_lookup_if_else_else_else_le_index_s_sva[5:0];
  assign _00453_ = _01127_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11589" *) _00857_ : lut_lookup_4_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  assign _00464_ = _01126_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11579" *) lut_lookup_else_1_lo_index_u_3_sva_3 : lut_lookup_else_1_lo_index_u_3_sva_4;
  assign _00508_ = _01125_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11571" *) lut_lookup_else_else_else_le_index_u_3_sva_3 : lut_lookup_else_else_else_le_index_u_3_sva_4;
  assign _00856_ = and_dcpl_148 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_else_else_else_lut_lookup_else_else_else_and_5_nl : lut_lookup_if_else_else_else_le_index_s_3_sva[5:0];
  assign _00427_ = _01124_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11561" *) _00856_ : lut_lookup_3_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  assign _00462_ = _01123_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11551" *) lut_lookup_else_1_lo_index_u_2_sva_3 : lut_lookup_else_1_lo_index_u_2_sva_4;
  assign _00506_ = _01122_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11543" *) lut_lookup_else_else_else_le_index_u_2_sva_3 : lut_lookup_else_else_else_le_index_u_2_sva_4;
  assign _00855_ = and_dcpl_148 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_else_else_else_lut_lookup_else_else_else_and_3_nl : lut_lookup_if_else_else_else_le_index_s_2_sva[5:0];
  assign _00402_ = _01121_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11533" *) _00855_ : lut_lookup_2_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  assign _00460_ = _01120_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11523" *) lut_lookup_else_1_lo_index_u_1_sva_3 : lut_lookup_else_1_lo_index_u_1_sva_4;
  assign _00504_ = _01119_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11515" *) lut_lookup_else_else_else_le_index_u_1_sva_3 : lut_lookup_else_else_else_le_index_u_1_sva_4;
  assign _00854_ = and_dcpl_148 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_else_else_else_lut_lookup_else_else_else_and_1_nl : lut_lookup_if_else_else_else_le_index_s_1_sva[5:0];
  assign _00377_ = _01118_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11505" *) _00854_ : lut_lookup_1_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2;
  assign _00256_ = IsNaN_8U_23U_8_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11494" *) IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_mx0w0 : IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_3_itm_2;
  assign _00265_ = IsNaN_8U_23U_8_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11494" *) IsNaN_8U_23U_8_nor_2_tmp_1 : IsNaN_8U_23U_8_nor_3_itm_2;
  assign _00777_ = and_dcpl_308 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _02146_ : chn_lut_in_rsci_d_mxwt[127];
  assign _00147_ = _01116_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11484" *) _00777_ : FpAdd_8U_23U_2_mux_49_itm_2;
  assign _00776_ = and_dcpl_316 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_mx0w0;
  assign _00222_ = _01115_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11475" *) _00776_ : IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2;
  assign _00228_ = _01114_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11466" *) IsNaN_8U_23U_4_nor_tmp : IsNaN_8U_23U_4_nor_3_itm_2;
  assign _00775_ = and_dcpl_304 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _02145_ : chn_lut_in_rsci_d_mxwt[127];
  assign _00115_ = _01113_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11457" *) _00775_ : FpAdd_8U_23U_1_mux_49_itm_2;
  assign _00255_ = IsNaN_8U_23U_8_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11448" *) IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_mx0w0 : IsNaN_8U_23U_8_IsNaN_8U_23U_8_nand_2_itm_2;
  assign _00264_ = IsNaN_8U_23U_8_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11448" *) IsNaN_8U_23U_8_nor_2_tmp_1 : IsNaN_8U_23U_8_nor_2_itm_2;
  assign _00774_ = and_dcpl_300 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _02146_ : chn_lut_in_rsci_d_mxwt[95];
  assign _00144_ = _01112_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11438" *) _00774_ : FpAdd_8U_23U_2_mux_33_itm_2;
  assign _00773_ = and_dcpl_296 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _02145_ : chn_lut_in_rsci_d_mxwt[95];
  assign _00112_ = _01111_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11429" *) _00773_ : FpAdd_8U_23U_1_mux_33_itm_2;
  assign _00772_ = and_dcpl_292 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _02146_ : chn_lut_in_rsci_d_mxwt[63];
  assign _00140_ = _01110_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11420" *) _00772_ : FpAdd_8U_23U_2_mux_17_itm_2;
  assign _00771_ = and_dcpl_288 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _02145_ : chn_lut_in_rsci_d_mxwt[63];
  assign _00108_ = _01108_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11411" *) _00771_ : FpAdd_8U_23U_1_mux_17_itm_2;
  assign _00770_ = and_dcpl_284 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _02146_ : chn_lut_in_rsci_d_mxwt[31];
  assign _00141_ = _01107_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11402" *) _00770_ : FpAdd_8U_23U_2_mux_1_itm_2;
  assign _00769_ = and_dcpl_316 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_mx0w0;
  assign _00223_ = _01106_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11393" *) _00769_ : IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2;
  assign _00229_ = _01104_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11384" *) IsNaN_8U_23U_4_nor_tmp : IsNaN_8U_23U_4_nor_itm_2;
  assign _00768_ = and_dcpl_280 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) _02145_ : chn_lut_in_rsci_d_mxwt[31];
  assign _00109_ = _01103_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11375" *) _00768_ : FpAdd_8U_23U_1_mux_1_itm_2;
  assign _00447_ = lut_lookup_lo_index_0_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11348" *) lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  assign _00421_ = lut_lookup_lo_index_0_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11348" *) lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  assign _00396_ = lut_lookup_lo_index_0_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11348" *) lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  assign _00371_ = lut_lookup_lo_index_0_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11348" *) lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3;
  assign _00626_ = lut_lookup_lo_index_0_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11348" *) _01101_ : lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_11;
  assign _00629_ = lut_lookup_lo_index_0_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11348" *) _01099_ : lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_11;
  assign _00632_ = lut_lookup_lo_index_0_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11348" *) _01097_ : lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_11;
  assign _00635_ = lut_lookup_lo_index_0_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11348" *) _01095_ : lut_lookup_lo_index_0_7_0_lpi_1_dfm_11;
  assign _00473_ = _01093_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11329" *) lut_lookup_else_1_slc_32_mdf_1_sva_6 : lut_lookup_else_1_slc_32_mdf_1_sva_7;
  assign _00477_ = lut_lookup_else_1_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11320" *) lut_lookup_else_1_slc_32_mdf_2_sva_6 : lut_lookup_else_1_slc_32_mdf_2_sva_7;
  assign _00481_ = lut_lookup_else_1_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11320" *) lut_lookup_else_1_slc_32_mdf_3_sva_6 : lut_lookup_else_1_slc_32_mdf_3_sva_7;
  assign _00485_ = _01092_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11311" *) lut_lookup_else_1_slc_32_mdf_sva_6 : lut_lookup_else_1_slc_32_mdf_sva_7;
  assign _00500_ = _01091_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11303" *) lut_lookup_4_else_else_else_if_acc_nl[3] : lut_lookup_else_else_else_asn_mdf_sva_3;
  assign _00193_ = _01090_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11295" *) lut_lookup_if_else_else_le_data_sub_sva_1_30_0_1 : IntLog2_32U_ac_int_cctor_1_30_0_sva_1;
  assign _00497_ = _01089_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11287" *) lut_lookup_3_else_else_else_if_acc_nl[3] : lut_lookup_else_else_else_asn_mdf_3_sva_3;
  assign _00192_ = _01088_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11279" *) lut_lookup_if_else_else_le_data_sub_3_sva_1_30_0_1 : IntLog2_32U_ac_int_cctor_1_30_0_3_sva_1;
  assign _00494_ = _01087_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11271" *) lut_lookup_2_else_else_else_if_acc_nl[3] : lut_lookup_else_else_else_asn_mdf_2_sva_3;
  assign _00517_ = lut_lookup_else_else_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11261" *) lut_lookup_2_if_else_slc_32_svs_6 : lut_lookup_else_else_slc_32_mdf_2_sva_7;
  assign _00519_ = lut_lookup_else_else_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11261" *) lut_lookup_3_if_else_slc_32_svs_6 : lut_lookup_else_else_slc_32_mdf_3_sva_7;
  assign _00521_ = lut_lookup_else_else_and_9_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11261" *) lut_lookup_4_if_else_slc_32_svs_6 : lut_lookup_else_else_slc_32_mdf_sva_7;
  assign _00191_ = _01086_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11251" *) lut_lookup_if_else_else_le_data_sub_2_sva_1_30_0_1 : IntLog2_32U_ac_int_cctor_1_30_0_2_sva_1;
  assign _00491_ = _01085_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11243" *) lut_lookup_1_else_else_else_if_acc_nl[3] : lut_lookup_else_else_else_asn_mdf_1_sva_3;
  assign _00515_ = _01084_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11235" *) lut_lookup_1_if_else_slc_32_svs_6 : lut_lookup_else_else_slc_32_mdf_1_sva_7;
  assign _00190_ = _01083_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11227" *) lut_lookup_if_else_else_le_data_sub_1_sva_1_30_0_1 : IntLog2_32U_ac_int_cctor_1_30_0_1_sva_2;
  assign _00767_ = and_679_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1 : _02140_;
  assign _00542_ = _01082_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11218" *) _00767_ : lut_lookup_else_mux_itm_2;
  assign _00766_ = and_428_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_if_lor_6_lpi_1_dfm_mx0w1 : _02139_;
  assign _00765_ = and_428_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_if_lor_7_lpi_1_dfm_mx0w1 : _02138_;
  assign _00764_ = and_428_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_if_lor_1_lpi_1_dfm_mx0w1 : _02137_;
  assign _00539_ = lut_lookup_else_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11205" *) _00764_ : lut_lookup_else_mux_129_itm_2;
  assign _00541_ = lut_lookup_else_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11205" *) _00765_ : lut_lookup_else_mux_86_itm_2;
  assign _00540_ = lut_lookup_else_and_8_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11205" *) _00766_ : lut_lookup_else_mux_43_itm_2;
  assign _00450_ = _01080_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11194" *) FpMantRNE_49U_24U_2_else_carry_sva_2 : lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign _00719_ = _01079_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11185" *) lut_lookup_else_1_else_else_mux1h_1_itm[7:0] : reg_lut_lookup_4_else_1_else_else_acc_1_itm;
  assign _00720_ = _01075_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11176" *) lut_lookup_else_1_else_else_mux1h_1_itm[8] : reg_lut_lookup_4_else_1_else_else_acc_itm;
  assign _00446_ = _01067_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11165" *) _01068_ : lut_lookup_4_else_1_else_else_lo_data_f_and_itm_2;
  assign _00849_ = and_676_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) FpAdd_8U_23U_2_asn_35_mx0w1 : lut_in_data_sva_156[118:96];
  assign _00157_ = _01066_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11156" *) _00849_ : FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5;
  assign _00501_ = _01063_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11147" *) lut_lookup_else_else_else_asn_mdf_sva_3 : lut_lookup_else_else_else_asn_mdf_sva_4;
  assign _00722_ = _01062_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11139" *) lut_lookup_else_else_else_else_mux1h_3_rgt[6:4] : reg_lut_lookup_4_else_else_else_else_acc_2_reg;
  assign _00451_ = _01059_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11129" *) _01060_ : lut_lookup_4_else_else_else_else_le_data_f_and_itm_2;
  assign _00444_ = _01058_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11120" *) reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[1:0] : lut_lookup_4_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  assign _00457_ = _01057_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11111" *) lut_lookup_4_if_else_slc_32_svs_7 : lut_lookup_4_if_else_slc_32_svs_8;
  assign _00580_ = _01056_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11103" *) lut_lookup_if_else_else_slc_10_mdf_sva_3 : lut_lookup_if_else_else_slc_10_mdf_sva_4;
  assign _00565_ = _01055_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11095" *) lut_lookup_4_if_else_else_else_if_acc_nl[3] : lut_lookup_if_else_else_else_asn_mdf_sva_2;
  assign _00582_ = _01054_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11087" *) lut_lookup_if_if_lor_1_lpi_1_dfm_mx0w3 : lut_lookup_if_if_lor_1_lpi_1_dfm_4;
  assign _00482_ = lut_lookup_else_1_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11078" *) lut_lookup_else_1_slc_32_mdf_3_sva_7 : lut_lookup_else_1_slc_32_mdf_3_sva_8;
  assign _00486_ = lut_lookup_else_1_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11078" *) lut_lookup_else_1_slc_32_mdf_sva_7 : lut_lookup_else_1_slc_32_mdf_sva_8;
  assign _00424_ = _01053_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11068" *) FpMantRNE_49U_24U_2_else_carry_3_sva_2 : lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign _00708_ = _01052_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11059" *) lut_lookup_else_1_else_else_mux1h_1_itm[7:0] : reg_lut_lookup_3_else_1_else_else_acc_1_itm;
  assign _00709_ = _01048_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11050" *) lut_lookup_else_1_else_else_mux1h_1_itm[8] : reg_lut_lookup_3_else_1_else_else_acc_itm;
  assign _00420_ = _01040_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11039" *) _01041_ : lut_lookup_3_else_1_else_else_lo_data_f_and_itm_2;
  assign _00848_ = and_668_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) FpAdd_8U_23U_2_asn_40_mx0w1 : lut_in_data_sva_156[86:64];
  assign _00156_ = _01039_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11030" *) _00848_ : FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5;
  assign _00498_ = _01036_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11021" *) lut_lookup_else_else_else_asn_mdf_3_sva_3 : lut_lookup_else_else_else_asn_mdf_3_sva_4;
  assign _00711_ = _01035_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11013" *) lut_lookup_else_else_else_else_mux1h_2_rgt[6:4] : reg_lut_lookup_3_else_else_else_else_acc_2_reg;
  assign _00425_ = _01032_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:11003" *) _01033_ : lut_lookup_3_else_else_else_else_le_data_f_and_itm_2;
  assign _00418_ = _01031_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10994" *) reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[1:0] : lut_lookup_3_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  assign _00577_ = _01030_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10985" *) lut_lookup_if_else_else_slc_10_mdf_3_sva_3 : lut_lookup_if_else_else_slc_10_mdf_3_sva_4;
  assign _00564_ = _01029_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10977" *) lut_lookup_3_if_else_else_else_if_acc_nl[3] : lut_lookup_if_else_else_else_asn_mdf_3_sva_2;
  assign _00478_ = _01028_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10969" *) lut_lookup_else_1_slc_32_mdf_2_sva_7 : lut_lookup_else_1_slc_32_mdf_2_sva_8;
  assign _00399_ = _01027_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10960" *) FpMantRNE_49U_24U_2_else_carry_2_sva_2 : lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign _00697_ = _01026_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10951" *) lut_lookup_else_1_else_else_mux1h_1_itm[7:0] : reg_lut_lookup_2_else_1_else_else_acc_1_itm;
  assign _00698_ = _01022_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10942" *) lut_lookup_else_1_else_else_mux1h_1_itm[8] : reg_lut_lookup_2_else_1_else_else_acc_itm;
  assign _00395_ = _01014_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10931" *) _01015_ : lut_lookup_2_else_1_else_else_lo_data_f_and_itm_2;
  assign _00847_ = and_661_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) FpAdd_8U_23U_2_asn_45_mx0w1 : lut_in_data_sva_156[54:32];
  assign _00155_ = _01013_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10922" *) _00847_ : FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5;
  assign _00518_ = lut_lookup_else_else_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10911" *) lut_lookup_else_else_slc_32_mdf_2_sva_7 : lut_lookup_else_else_slc_32_mdf_2_sva_8;
  assign _00520_ = lut_lookup_else_else_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10911" *) lut_lookup_else_else_slc_32_mdf_3_sva_7 : lut_lookup_else_else_slc_32_mdf_3_sva_8;
  assign _00522_ = lut_lookup_else_else_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10911" *) lut_lookup_else_else_slc_32_mdf_sva_7 : lut_lookup_else_else_slc_32_mdf_sva_8;
  assign _00495_ = _01010_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10901" *) lut_lookup_else_else_else_asn_mdf_2_sva_3 : lut_lookup_else_else_else_asn_mdf_2_sva_4;
  assign _00700_ = _01009_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10893" *) lut_lookup_else_else_else_else_mux1h_1_rgt[6:4] : reg_lut_lookup_2_else_else_else_else_acc_2_reg;
  assign _00400_ = _01006_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10883" *) { _02027_[31:6], _01007_ } : lut_lookup_2_else_else_else_else_le_data_f_and_itm_2;
  assign _00393_ = _01005_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10874" *) reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[1:0] : lut_lookup_2_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  assign _00675_ = and_907_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10863" *) IntLog2_32U_IntLog2_32U_mux_2_rgt[30:23] : reg_IntLog2_32U_ac_int_cctor_1_30_0_reg;
  assign _00674_ = and_907_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10863" *) IntLog2_32U_IntLog2_32U_mux_1_rgt[30:23] : reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg;
  assign _00671_ = and_907_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10863" *) IntLog2_32U_IntLog2_32U_mux_rgt[30:23] : reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg;
  assign _00574_ = _01004_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10853" *) lut_lookup_if_else_else_slc_10_mdf_2_sva_3 : lut_lookup_if_else_else_slc_10_mdf_2_sva_4;
  assign _00563_ = _01003_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10845" *) lut_lookup_2_if_else_else_else_if_acc_nl[3] : lut_lookup_if_else_else_else_asn_mdf_2_sva_2;
  assign _00474_ = _01002_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10837" *) lut_lookup_else_1_slc_32_mdf_1_sva_7 : lut_lookup_else_1_slc_32_mdf_1_sva_8;
  assign _00374_ = _01001_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10828" *) FpMantRNE_49U_24U_2_else_carry_1_sva_2 : lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_4_itm_3;
  assign _00686_ = _01000_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10819" *) lut_lookup_else_1_else_else_mux1h_1_itm[7:0] : reg_lut_lookup_1_else_1_else_else_acc_1_itm;
  assign _00687_ = _00996_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10810" *) lut_lookup_else_1_else_else_mux1h_1_itm[8] : reg_lut_lookup_1_else_1_else_else_acc_itm;
  assign _00370_ = _00988_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10799" *) _00989_ : lut_lookup_1_else_1_else_else_lo_data_f_and_itm_2;
  assign _00846_ = and_653_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13493|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13492" *) FpAdd_8U_23U_2_asn_50_mx0w1 : lut_in_data_sva_156[22:0];
  assign _00154_ = _00987_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10790" *) _00846_ : FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5;
  assign _00516_ = _00984_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10781" *) lut_lookup_else_else_slc_32_mdf_1_sva_7 : lut_lookup_else_else_slc_32_mdf_1_sva_8;
  assign _00492_ = _00983_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10773" *) lut_lookup_else_else_else_asn_mdf_1_sva_3 : lut_lookup_else_else_else_asn_mdf_1_sva_4;
  assign _00723_ = and_905_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10759" *) lut_lookup_else_else_else_else_mux1h_3_rgt[3:0] : reg_lut_lookup_4_else_else_else_else_acc_3_reg;
  assign _00672_ = and_905_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10759" *) IntLog2_32U_IntLog2_32U_mux_2_rgt[22:0] : reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1;
  assign _00712_ = and_905_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10759" *) lut_lookup_else_else_else_else_mux1h_2_rgt[3:0] : reg_lut_lookup_3_else_else_else_else_acc_3_reg;
  assign _00673_ = and_905_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10759" *) IntLog2_32U_IntLog2_32U_mux_1_rgt[22:0] : reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg;
  assign _00701_ = and_905_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10759" *) lut_lookup_else_else_else_else_mux1h_1_rgt[3:0] : reg_lut_lookup_2_else_else_else_else_acc_3_reg;
  assign _00670_ = and_905_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10759" *) IntLog2_32U_IntLog2_32U_mux_rgt[22:0] : reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg;
  assign _00690_ = and_905_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10759" *) lut_lookup_else_else_else_else_mux1h_rgt[3:0] : reg_lut_lookup_1_else_else_else_else_acc_3_reg;
  assign _00689_ = _00982_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10745" *) lut_lookup_else_else_else_else_mux1h_rgt[6:4] : reg_lut_lookup_1_else_else_else_else_acc_2_reg;
  assign _00721_ = and_901_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10733" *) lut_lookup_else_else_else_else_mux1h_3_rgt[7] : reg_lut_lookup_4_else_else_else_else_acc_1_reg;
  assign _00710_ = and_901_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10733" *) lut_lookup_else_else_else_else_mux1h_2_rgt[7] : reg_lut_lookup_3_else_else_else_else_acc_1_reg;
  assign _00699_ = and_901_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10733" *) lut_lookup_else_else_else_else_mux1h_1_rgt[7] : reg_lut_lookup_2_else_else_else_else_acc_1_reg;
  assign _00688_ = and_901_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10733" *) lut_lookup_else_else_else_else_mux1h_rgt[7] : reg_lut_lookup_1_else_else_else_else_acc_1_reg;
  assign _00724_ = and_898_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10719" *) lut_lookup_else_else_else_else_mux1h_3_rgt[8] : reg_lut_lookup_4_else_else_else_else_acc_reg;
  assign _00713_ = and_898_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10719" *) lut_lookup_else_else_else_else_mux1h_2_rgt[8] : reg_lut_lookup_3_else_else_else_else_acc_reg;
  assign _00702_ = and_898_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10719" *) lut_lookup_else_else_else_else_mux1h_1_rgt[8] : reg_lut_lookup_2_else_else_else_else_acc_reg;
  assign _00691_ = and_898_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10719" *) lut_lookup_else_else_else_else_mux1h_rgt[8] : reg_lut_lookup_1_else_else_else_else_acc_reg;
  assign _00375_ = _00979_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10707" *) _00980_ : lut_lookup_1_else_else_else_else_le_data_f_and_itm_2;
  assign _00300_ = _00978_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10699" *) cfg_precision_1_sva_st_70 : cfg_precision_1_sva_8;
  assign _00368_ = _00977_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10690" *) reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[1:0] : lut_lookup_1_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3;
  assign _00668_ = _00976_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10681" *) IntLog2_32U_mux1h_1_itm[22:0] : reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm;
  assign _00669_ = _00974_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10673" *) IntLog2_32U_mux1h_1_itm[30:23] : reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm;
  assign _00381_ = lut_lookup_if_else_if_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10660" *) lut_lookup_1_if_else_slc_32_svs_7 : lut_lookup_1_if_else_slc_32_svs_8;
  assign _00406_ = lut_lookup_if_else_if_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10660" *) lut_lookup_2_if_else_slc_32_svs_7 : lut_lookup_2_if_else_slc_32_svs_8;
  assign _00431_ = lut_lookup_if_else_if_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10660" *) lut_lookup_3_if_else_slc_32_svs_7 : lut_lookup_3_if_else_slc_32_svs_8;
  assign _00571_ = _00967_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10650" *) lut_lookup_if_else_else_slc_10_mdf_1_sva_3 : lut_lookup_if_else_else_slc_10_mdf_1_sva_4;
  assign _00562_ = _00966_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10642" *) lut_lookup_1_if_else_else_else_if_acc_nl[3] : lut_lookup_if_else_else_else_asn_mdf_1_sva_2;
  assign _00583_ = lut_lookup_if_if_oelse_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10632" *) lut_lookup_if_if_lor_5_lpi_1_dfm_mx0w3 : lut_lookup_if_if_lor_5_lpi_1_dfm_4;
  assign _00584_ = lut_lookup_if_if_oelse_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10632" *) lut_lookup_if_if_lor_6_lpi_1_dfm_mx0w3 : lut_lookup_if_if_lor_6_lpi_1_dfm_4;
  assign _00585_ = lut_lookup_if_if_oelse_1_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10632" *) lut_lookup_if_if_lor_7_lpi_1_dfm_mx0w3 : lut_lookup_if_if_lor_7_lpi_1_dfm_4;
  assign _00763_ = and_427_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5 : and_1141_cse;
  assign _00194_ = _00965_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10621" *) _00763_ : IsNaN_8U_23U_10_land_1_lpi_1_dfm_5;
  assign _00553_ = lut_lookup_if_1_oelse_1_and_14_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10611" *) or_969_cse : lut_lookup_if_1_lor_5_lpi_1_dfm_4;
  assign _00556_ = lut_lookup_if_1_oelse_1_and_14_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10611" *) lut_lookup_if_1_lor_6_lpi_1_dfm_mx0w0 : lut_lookup_if_1_lor_6_lpi_1_dfm_4;
  assign _00762_ = and_427_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5 : and_1140_cse;
  assign _00196_ = _00964_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10601" *) _00762_ : IsNaN_8U_23U_10_land_2_lpi_1_dfm_5;
  assign _00397_ = lut_lookup_lo_index_0_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10587" *) lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 : lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  assign _00372_ = lut_lookup_lo_index_0_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10587" *) lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 : lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  assign _00627_ = lut_lookup_lo_index_0_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10587" *) lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_11 : lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_12;
  assign _00630_ = lut_lookup_lo_index_0_and_6_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10587" *) lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_11 : lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_12;
  assign _00761_ = and_427_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5 : and_1139_cse;
  assign _00198_ = _00963_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10573" *) _00761_ : IsNaN_8U_23U_10_land_3_lpi_1_dfm_5;
  assign _00559_ = lut_lookup_if_1_oelse_1_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10563" *) lut_lookup_if_1_lor_7_lpi_1_dfm_mx0w0 : lut_lookup_if_1_lor_7_lpi_1_dfm_4;
  assign _00550_ = lut_lookup_if_1_oelse_1_and_12_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10563" *) lut_lookup_if_1_lor_1_lpi_1_dfm_mx0w0 : lut_lookup_if_1_lor_1_lpi_1_dfm_4;
  assign _00760_ = and_427_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5 : and_1138_cse;
  assign _00200_ = _00962_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10553" *) _00760_ : IsNaN_8U_23U_10_land_lpi_1_dfm_5;
  assign _00448_ = lut_lookup_lo_index_0_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10539" *) lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 : lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  assign _00422_ = lut_lookup_lo_index_0_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10539" *) lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_3 : lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_1_itm_4;
  assign _00633_ = lut_lookup_lo_index_0_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10539" *) lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_11 : lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_12;
  assign _00636_ = lut_lookup_lo_index_0_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10539" *) lut_lookup_lo_index_0_7_0_lpi_1_dfm_11 : lut_lookup_lo_index_0_7_0_lpi_1_dfm_12;
  assign _00530_ = _00960_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10526" *) lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1 : lut_lookup_else_if_lor_5_lpi_1_dfm_5;
  assign _00230_ = _00959_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10516" *) _03226_ : IsNaN_8U_23U_6_land_1_lpi_1_dfm_6;
  assign _00232_ = _00958_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10504" *) _03225_ : IsNaN_8U_23U_6_land_2_lpi_1_dfm_6;
  assign _00234_ = _00957_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10492" *) _03224_ : IsNaN_8U_23U_6_land_3_lpi_1_dfm_6;
  assign _00543_ = _00956_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10483" *) lut_lookup_unequal_tmp_mx0w0 : lut_lookup_else_unequal_tmp_12;
  assign _00533_ = lut_lookup_else_if_oelse_1_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10473" *) lut_lookup_else_if_lor_6_lpi_1_dfm_mx0w1 : lut_lookup_else_if_lor_6_lpi_1_dfm_5;
  assign _00536_ = lut_lookup_else_if_oelse_1_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10473" *) lut_lookup_else_if_lor_7_lpi_1_dfm_mx0w1 : lut_lookup_else_if_lor_7_lpi_1_dfm_5;
  assign _00527_ = lut_lookup_else_if_oelse_1_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10473" *) lut_lookup_else_if_lor_1_lpi_1_dfm_mx0w1 : lut_lookup_else_if_lor_1_lpi_1_dfm_5;
  assign _00236_ = _00955_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10460" *) _03223_ : IsNaN_8U_23U_6_land_lpi_1_dfm_6;
  assign _00465_ = _00953_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10451" *) nl_lut_lookup_else_1_lo_index_u_sva_3[31:0] : lut_lookup_else_1_lo_index_u_sva_3;
  assign _00509_ = _00952_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10443" *) lut_lookup_if_else_else_le_data_sub_sva_mx0w0 : lut_lookup_else_else_else_le_index_u_sva_3;
  assign _00463_ = _00951_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10435" *) nl_lut_lookup_else_1_lo_index_u_3_sva_3[31:0] : lut_lookup_else_1_lo_index_u_3_sva_3;
  assign _00507_ = _00950_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10427" *) lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0 : lut_lookup_else_else_else_le_index_u_3_sva_3;
  assign _00461_ = _00949_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10419" *) nl_lut_lookup_else_1_lo_index_u_2_sva_3 : lut_lookup_else_1_lo_index_u_2_sva_3;
  assign _00505_ = _00948_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10411" *) lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0 : lut_lookup_else_else_else_le_index_u_2_sva_3;
  assign _00459_ = _00947_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10403" *) nl_lut_lookup_else_1_lo_index_u_1_sva_3 : lut_lookup_else_1_lo_index_u_1_sva_3;
  assign _00503_ = _00946_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10395" *) lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0 : lut_lookup_else_else_else_le_index_u_1_sva_3;
  assign _00148_ = _00945_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10385" *) _03222_ : FpAdd_8U_23U_2_mux_61_itm_1;
  assign _00116_ = _00943_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10374" *) _03202_ : FpAdd_8U_23U_1_mux_61_itm_3;
  assign _00145_ = _00941_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10363" *) _03221_ : FpAdd_8U_23U_2_mux_45_itm_1;
  assign _00113_ = _00939_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10352" *) _03201_ : FpAdd_8U_23U_1_mux_45_itm_3;
  assign _00142_ = _00937_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10341" *) _03220_ : FpAdd_8U_23U_2_mux_29_itm_1;
  assign _00110_ = _00935_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10330" *) _03200_ : FpAdd_8U_23U_1_mux_29_itm_3;
  assign _00138_ = _00933_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10319" *) _03219_ : FpAdd_8U_23U_2_mux_13_itm_1;
  assign _00106_ = _00931_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10308" *) _03199_ : FpAdd_8U_23U_1_mux_13_itm_3;
  assign _00759_ = and_525_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4 : reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse;
  assign _00758_ = and_525_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4 : IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  assign _00757_ = and_525_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4 : IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
  assign _00252_ = IsNaN_8U_23U_1_aelse_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10294" *) _00759_ : IsNaN_8U_23U_7_land_lpi_1_dfm_6;
  assign _00247_ = IsNaN_8U_23U_1_aelse_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10294" *) _00758_ : IsNaN_8U_23U_7_land_3_lpi_1_dfm_6;
  assign _00243_ = IsNaN_8U_23U_1_aelse_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10294" *) _00757_ : IsNaN_8U_23U_7_land_2_lpi_1_dfm_6;
  assign _00756_ = and_524_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_itm_2 : IsNaN_8U_23U_4_land_1_lpi_1_dfm_mx0w0;
  assign _00224_ = _00929_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10283" *) _00756_ : IsNaN_8U_23U_4_land_1_lpi_1_dfm_4;
  assign _00206_ = IsNaN_8U_23U_1_aelse_and_5_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10269" *) _03198_ : IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _00208_ = IsNaN_8U_23U_1_aelse_and_5_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10269" *) _03197_ : IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign _00755_ = and_525_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4 : IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
  assign _00754_ = and_525_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 : IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _00753_ = and_525_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 : IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _00238_ = IsNaN_8U_23U_1_aelse_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10255" *) _00755_ : IsNaN_8U_23U_7_land_1_lpi_1_dfm_6;
  assign _00203_ = IsNaN_8U_23U_1_aelse_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10255" *) _00754_ : IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign _00211_ = IsNaN_8U_23U_1_aelse_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10255" *) _00753_ : IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _00752_ = and_524_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4 : IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _00751_ = and_524_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4 : IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _00750_ = and_524_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_3_itm_2 : IsNaN_8U_23U_4_land_lpi_1_dfm_mx0w0;
  assign _00225_ = IsNaN_8U_23U_3_aelse_and_3_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10240" *) _00752_ : IsNaN_8U_23U_4_land_2_lpi_1_dfm_5;
  assign _00226_ = IsNaN_8U_23U_3_aelse_and_3_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10240" *) _00751_ : IsNaN_8U_23U_4_land_3_lpi_1_dfm_5;
  assign _00227_ = IsNaN_8U_23U_3_aelse_and_3_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10240" *) _00750_ : IsNaN_8U_23U_4_land_lpi_1_dfm_4;
  assign _00125_ = _00927_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10230" *) acc_5_nl[8:1] : FpAdd_8U_23U_2_a_right_shift_qr_sva_3;
  assign _00436_ = IsZero_8U_23U_7_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10221" *) _02055_ : lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2;
  assign _00435_ = IsZero_8U_23U_7_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10221" *) lut_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 : lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  assign _00124_ = _00926_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10212" *) acc_9_nl[8:1] : FpAdd_8U_23U_2_a_right_shift_qr_3_sva_3;
  assign _00410_ = _00925_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10204" *) lut_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 : lut_lookup_3_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  assign _00749_ = and_dcpl_315 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
  assign _00748_ = and_dcpl_316 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 : lut_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  assign _00747_ = and_dcpl_316 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 : lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  assign _00746_ = and_dcpl_316 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 : lut_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  assign _00745_ = and_dcpl_316 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 : lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  assign _00744_ = and_dcpl_316 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 : lut_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  assign _00743_ = and_dcpl_316 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 : lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  assign _00434_ = IsZero_8U_23U_4_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10183" *) _00747_ : lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  assign _00433_ = IsZero_8U_23U_4_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10183" *) _00748_ : lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  assign _00409_ = IsZero_8U_23U_4_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10183" *) _00745_ : lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  assign _00408_ = IsZero_8U_23U_4_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10183" *) _00746_ : lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  assign _00384_ = IsZero_8U_23U_4_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10183" *) _00743_ : lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  assign _00383_ = IsZero_8U_23U_4_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10183" *) _00744_ : lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  assign _00210_ = IsZero_8U_23U_4_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10183" *) _00749_ : IsNaN_8U_23U_1_land_lpi_1_dfm_6;
  assign _00742_ = and_dcpl_314 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_4_else_1_acc_nl[32] : FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_3_cse;
  assign _00741_ = and_dcpl_314 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_3_else_1_acc_nl[32] : FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_2_cse;
  assign _00740_ = and_dcpl_314 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_2_else_1_acc_nl[32] : FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_1_cse;
  assign _00739_ = and_dcpl_314 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_1_else_1_acc_nl[32] : FpAdd_8U_23U_2_is_a_greater_FpAdd_8U_23U_2_is_a_greater_or_cse;
  assign _00133_ = FpAdd_8U_23U_2_is_a_greater_oelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10162" *) _00742_ : FpAdd_8U_23U_2_is_a_greater_lor_lpi_1_dfm_4;
  assign _00132_ = FpAdd_8U_23U_2_is_a_greater_oelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10162" *) _00741_ : FpAdd_8U_23U_2_is_a_greater_lor_3_lpi_1_dfm_4;
  assign _00131_ = FpAdd_8U_23U_2_is_a_greater_oelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10162" *) _00740_ : FpAdd_8U_23U_2_is_a_greater_lor_2_lpi_1_dfm_4;
  assign _00130_ = FpAdd_8U_23U_2_is_a_greater_oelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10162" *) _00739_ : FpAdd_8U_23U_2_is_a_greater_lor_1_lpi_1_dfm_4;
  assign _00738_ = and_dcpl_315 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0;
  assign _00737_ = and_dcpl_316 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0 : lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1;
  assign _00736_ = and_dcpl_316 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 : lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_mx0w0;
  assign _00359_ = IsZero_8U_23U_4_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10146" *) _00736_ : lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2;
  assign _00358_ = IsZero_8U_23U_4_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10146" *) _00737_ : lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  assign _00202_ = IsZero_8U_23U_4_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10146" *) _00738_ : IsNaN_8U_23U_1_land_1_lpi_1_dfm_6;
  assign _00735_ = and_dcpl_314 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_4_else_else_acc_1_nl[32] : FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_3_cse;
  assign _00734_ = and_dcpl_314 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_3_else_else_acc_1_nl[32] : FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_2_cse;
  assign _00733_ = and_dcpl_314 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_2_else_else_acc_1_nl[32] : FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_1_cse;
  assign _00732_ = and_dcpl_314 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_1_else_else_acc_1_nl[32] : FpAdd_8U_23U_1_is_a_greater_FpAdd_8U_23U_1_is_a_greater_or_cse;
  assign _00101_ = FpAdd_8U_23U_1_is_a_greater_oelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10129" *) _00735_ : FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5;
  assign _00100_ = FpAdd_8U_23U_1_is_a_greater_oelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10129" *) _00734_ : FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5;
  assign _00099_ = FpAdd_8U_23U_1_is_a_greater_oelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10129" *) _00733_ : FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5;
  assign _00098_ = FpAdd_8U_23U_1_is_a_greater_oelse_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10129" *) _00732_ : FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5;
  assign _00865_ = and_dcpl_308 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) cfg_lut_lo_start_rsci_d[30:23] : chn_lut_in_rsci_d_mxwt[126:119];
  assign _00164_ = _00923_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10117" *) _00865_ : FpAdd_8U_23U_2_qr_lpi_1_dfm_4;
  assign _00864_ = and_dcpl_300 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) cfg_lut_lo_start_rsci_d[30:23] : chn_lut_in_rsci_d_mxwt[94:87];
  assign _00162_ = _00921_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10108" *) _00864_ : FpAdd_8U_23U_2_qr_4_lpi_1_dfm_4;
  assign _00863_ = and_dcpl_292 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) cfg_lut_lo_start_rsci_d[30:23] : chn_lut_in_rsci_d_mxwt[62:55];
  assign _00160_ = FpAdd_8U_23U_2_and_44_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10098" *) _00863_ : FpAdd_8U_23U_2_qr_3_lpi_1_dfm_4;
  assign _00123_ = FpAdd_8U_23U_2_and_44_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10098" *) acc_10_nl[8:1] : FpAdd_8U_23U_2_a_right_shift_qr_2_sva_3;
  assign _00862_ = and_dcpl_280 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) cfg_lut_le_start_rsci_d[30:23] : chn_lut_in_rsci_d_mxwt[30:23];
  assign _00118_ = FpAdd_8U_23U_1_and_46_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10087" *) _00862_ : FpAdd_8U_23U_1_qr_2_lpi_1_dfm_5;
  assign _00090_ = FpAdd_8U_23U_1_and_46_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10087" *) acc_4_nl[8:1] : FpAdd_8U_23U_1_a_right_shift_qr_1_sva_3;
  assign _00731_ = and_428_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_1_lor_1_lpi_1_dfm_mx0w0 : _02099_;
  assign _00730_ = and_428_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_1_lor_7_lpi_1_dfm_mx0w0 : _02098_;
  assign _00729_ = and_428_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_1_lor_6_lpi_1_dfm_mx0w0 : _02097_;
  assign _00728_ = and_428_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) or_969_cse : _02096_;
  assign _00644_ = lut_lookup_lo_uflow_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10071" *) _00731_ : lut_lookup_lo_uflow_lpi_1_dfm_3;
  assign _00642_ = lut_lookup_lo_uflow_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10071" *) _00730_ : lut_lookup_lo_uflow_3_lpi_1_dfm_3;
  assign _00640_ = lut_lookup_lo_uflow_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10071" *) _00729_ : lut_lookup_lo_uflow_2_lpi_1_dfm_3;
  assign _00638_ = lut_lookup_lo_uflow_and_4_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10071" *) _00728_ : lut_lookup_lo_uflow_1_lpi_1_dfm_3;
  assign _00512_ = _00919_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10058" *) _03196_ : lut_lookup_else_else_lut_lookup_else_else_and_1_itm_2;
  assign _00469_ = lut_lookup_lo_index_0_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10044" *) _00916_ : lut_lookup_else_1_lut_lookup_else_1_and_4_itm_2;
  assign _00468_ = lut_lookup_lo_index_0_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10044" *) _00917_ : lut_lookup_else_1_lut_lookup_else_1_and_1_itm_2;
  assign _00628_ = lut_lookup_lo_index_0_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10044" *) lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_12 : lut_lookup_lo_index_0_7_0_1_lpi_1_dfm_13;
  assign _00631_ = lut_lookup_lo_index_0_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10044" *) lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_12 : lut_lookup_lo_index_0_7_0_2_lpi_1_dfm_13;
  assign _00511_ = lut_lookup_else_else_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10025" *) _03193_ : lut_lookup_else_else_lut_lookup_else_else_and_10_itm_2;
  assign _00514_ = lut_lookup_else_else_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10025" *) _03194_ : lut_lookup_else_else_lut_lookup_else_else_and_7_itm_2;
  assign _00513_ = lut_lookup_else_else_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10025" *) _03195_ : lut_lookup_else_else_lut_lookup_else_else_and_4_itm_2;
  assign _00467_ = lut_lookup_lo_index_0_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10010" *) _00914_ : lut_lookup_else_1_lut_lookup_else_1_and_10_itm_2;
  assign _00470_ = lut_lookup_lo_index_0_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10010" *) _00915_ : lut_lookup_else_1_lut_lookup_else_1_and_7_itm_2;
  assign _00634_ = lut_lookup_lo_index_0_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10010" *) lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_12 : lut_lookup_lo_index_0_7_0_3_lpi_1_dfm_13;
  assign _00637_ = lut_lookup_lo_index_0_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:10010" *) lut_lookup_lo_index_0_7_0_lpi_1_dfm_12 : lut_lookup_lo_index_0_7_0_lpi_1_dfm_13;
  assign _00841_ = and_dcpl_259 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_mux_mx0w1 : lut_lookup_else_mux_itm_2;
  assign _00840_ = and_dcpl_259 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_mux_41_mx0w1 : lut_lookup_else_mux_43_itm_2;
  assign _00839_ = and_dcpl_259 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_mux_82_mx0w1 : lut_lookup_else_mux_86_itm_2;
  assign _00838_ = and_dcpl_259 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_if_mux_123_mx0w1 : lut_lookup_else_mux_129_itm_2;
  assign _00621_ = lut_lookup_le_uflow_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9992" *) _00838_ : lut_lookup_le_uflow_lpi_1_dfm_6;
  assign _00620_ = lut_lookup_le_uflow_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9992" *) _00839_ : lut_lookup_le_uflow_3_lpi_1_dfm_6;
  assign _00619_ = lut_lookup_le_uflow_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9992" *) _00840_ : lut_lookup_le_uflow_2_lpi_1_dfm_6;
  assign _00618_ = lut_lookup_le_uflow_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9992" *) _00841_ : lut_lookup_le_uflow_1_lpi_1_dfm_6;
  assign _00173_ = _02026_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9981" *) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_sva_2;
  assign _00201_ = _02025_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9973" *) IsNaN_8U_23U_10_land_lpi_1_dfm_5 : IsNaN_8U_23U_10_land_lpi_1_dfm_6;
  assign _00438_ = _02024_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9964" *) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9] : lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  assign _00549_ = _02023_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9955" *) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm : lut_lookup_if_1_else_lo_fra_sva_4;
  assign _00181_ = _02022_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9947" *) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm : FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_sva_2;
  assign _00237_ = _02021_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9939" *) IsNaN_8U_23U_6_land_lpi_1_dfm_6 : IsNaN_8U_23U_6_land_lpi_1_dfm_7;
  assign _00440_ = _02020_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9930" *) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9] : lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  assign _00526_ = _02019_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9921" *) lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm : lut_lookup_else_if_else_le_fra_sva_4;
  assign _00837_ = lut_lookup_else_2_else_else_if_mux_26_itm_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_186_cse : lut_lookup_lo_uflow_lpi_1_dfm_3;
  assign _00489_ = _02018_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9912" *) _00837_ : lut_lookup_else_2_else_else_if_mux_26_itm_1;
  assign _00560_ = lut_lookup_if_1_oelse_1_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9902" *) lut_lookup_if_1_lor_7_lpi_1_dfm_4 : lut_lookup_if_1_lor_7_lpi_1_dfm_5;
  assign _00551_ = lut_lookup_if_1_oelse_1_and_8_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9902" *) lut_lookup_if_1_lor_1_lpi_1_dfm_4 : lut_lookup_if_1_lor_1_lpi_1_dfm_5;
  assign _00172_ = _02016_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9893" *) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_3_sva_2;
  assign _00199_ = _02015_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9885" *) IsNaN_8U_23U_10_land_3_lpi_1_dfm_5 : IsNaN_8U_23U_10_land_3_lpi_1_dfm_6;
  assign _00412_ = _02014_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9876" *) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9] : lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  assign _00548_ = _02013_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9867" *) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm : lut_lookup_if_1_else_lo_fra_3_sva_4;
  assign _00537_ = lut_lookup_else_if_oelse_1_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9858" *) lut_lookup_else_if_lor_7_lpi_1_dfm_5 : lut_lookup_else_if_lor_7_lpi_1_dfm_6;
  assign _00528_ = lut_lookup_else_if_oelse_1_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9858" *) lut_lookup_else_if_lor_1_lpi_1_dfm_5 : lut_lookup_else_if_lor_1_lpi_1_dfm_6;
  assign _00180_ = _02012_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9849" *) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm : FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_3_sva_2;
  assign _00235_ = _02011_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9841" *) IsNaN_8U_23U_6_land_3_lpi_1_dfm_6 : IsNaN_8U_23U_6_land_3_lpi_1_dfm_7;
  assign _00414_ = _02010_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9832" *) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9] : lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  assign _00525_ = _02009_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9823" *) lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm : lut_lookup_else_if_else_le_fra_3_sva_4;
  assign _00836_ = lut_lookup_else_2_else_else_if_mux_19_itm_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_184_cse : lut_lookup_lo_uflow_3_lpi_1_dfm_3;
  assign _00488_ = _02008_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9814" *) _00836_ : lut_lookup_else_2_else_else_if_mux_19_itm_1;
  assign _00171_ = _02006_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9805" *) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_2_sva_2;
  assign _00197_ = _02005_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9797" *) IsNaN_8U_23U_10_land_2_lpi_1_dfm_5 : IsNaN_8U_23U_10_land_2_lpi_1_dfm_6;
  assign _00387_ = _02004_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9788" *) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9] : lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  assign _00547_ = _02003_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9779" *) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm : lut_lookup_if_1_else_lo_fra_2_sva_4;
  assign _00535_ = _02002_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9771" *) lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 : lut_lookup_else_if_lor_6_lpi_1_dfm_st_3;
  assign _00534_ = _02001_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9763" *) lut_lookup_else_if_lor_6_lpi_1_dfm_5 : lut_lookup_else_if_lor_6_lpi_1_dfm_6;
  assign _00179_ = _02000_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9755" *) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm : FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_2_sva_2;
  assign _00233_ = _01999_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9747" *) IsNaN_8U_23U_6_land_2_lpi_1_dfm_6 : IsNaN_8U_23U_6_land_2_lpi_1_dfm_7;
  assign _00389_ = _01998_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9738" *) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9] : lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  assign _00524_ = _01997_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9729" *) lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm : lut_lookup_else_if_else_le_fra_2_sva_4;
  assign _00835_ = lut_lookup_else_2_else_else_if_mux_12_itm_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_182_cse : lut_lookup_lo_uflow_2_lpi_1_dfm_3;
  assign _00487_ = _01996_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9720" *) _00835_ : lut_lookup_else_2_else_else_if_mux_12_itm_1;
  assign _00552_ = lut_lookup_if_1_oelse_1_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9708" *) lut_lookup_if_1_lor_1_lpi_1_dfm_4 : lut_lookup_if_1_lor_1_lpi_1_dfm_st_4;
  assign _00561_ = lut_lookup_if_1_oelse_1_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9708" *) lut_lookup_if_1_lor_7_lpi_1_dfm_4 : lut_lookup_if_1_lor_7_lpi_1_dfm_st_4;
  assign _00558_ = lut_lookup_if_1_oelse_1_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9708" *) lut_lookup_if_1_lor_6_lpi_1_dfm_4 : lut_lookup_if_1_lor_6_lpi_1_dfm_st_4;
  assign _00555_ = lut_lookup_if_1_oelse_1_and_5_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9708" *) lut_lookup_if_1_lor_5_lpi_1_dfm_4 : lut_lookup_if_1_lor_5_lpi_1_dfm_st_4;
  assign _00554_ = lut_lookup_if_1_oelse_1_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9696" *) lut_lookup_if_1_lor_5_lpi_1_dfm_4 : lut_lookup_if_1_lor_5_lpi_1_dfm_5;
  assign _00557_ = lut_lookup_if_1_oelse_1_and_4_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9696" *) lut_lookup_if_1_lor_6_lpi_1_dfm_4 : lut_lookup_if_1_lor_6_lpi_1_dfm_5;
  assign _00170_ = _01994_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9687" *) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_1_sva_2;
  assign _00195_ = _01993_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9679" *) IsNaN_8U_23U_10_land_1_lpi_1_dfm_5 : IsNaN_8U_23U_10_land_1_lpi_1_dfm_6;
  assign _00362_ = _01992_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9670" *) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9] : lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_9_itm_2;
  assign _00546_ = _01991_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9661" *) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm : lut_lookup_if_1_else_lo_fra_1_sva_4;
  assign _00304_ = _01990_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9653" *) cfg_precision_1_sva_st_71 : cfg_precision_1_sva_st_72;
  assign _00529_ = lut_lookup_else_if_oelse_1_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9643" *) lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 : lut_lookup_else_if_lor_1_lpi_1_dfm_st_3;
  assign _00538_ = lut_lookup_else_if_oelse_1_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9643" *) lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 : lut_lookup_else_if_lor_7_lpi_1_dfm_st_3;
  assign _00532_ = lut_lookup_else_if_oelse_1_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9643" *) lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2 : lut_lookup_else_if_lor_5_lpi_1_dfm_st_3;
  assign _00531_ = _01989_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9633" *) lut_lookup_else_if_lor_5_lpi_1_dfm_5 : lut_lookup_else_if_lor_5_lpi_1_dfm_6;
  assign _00178_ = _01988_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9625" *) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm : FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_1_sva_2;
  assign _00231_ = _01987_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9617" *) IsNaN_8U_23U_6_land_1_lpi_1_dfm_6 : IsNaN_8U_23U_6_land_1_lpi_1_dfm_7;
  assign _00364_ = _01986_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9608" *) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9] : lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_slc_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_9_itm_2;
  assign _00523_ = _01985_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9599" *) lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm : lut_lookup_else_if_else_le_fra_1_sva_4;
  assign _00834_ = lut_lookup_else_2_else_else_if_mux_5_itm_1_mx0c1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_mux_180_cse : lut_lookup_lo_uflow_1_lpi_1_dfm_3;
  assign _00490_ = _01984_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9590" *) _00834_ : lut_lookup_else_2_else_else_if_mux_5_itm_1;
  assign _00727_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_if_unequal_tmp_1_mx0w0 : reg_lut_lookup_if_unequal_cse;
  assign _00586_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01929_ : lut_lookup_le_fraction_1_lpi_1_dfm_16_34_12_1;
  assign _00589_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01939_ : lut_lookup_le_fraction_2_lpi_1_dfm_16_34_12_1;
  assign _00592_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01949_ : lut_lookup_le_fraction_3_lpi_1_dfm_16_34_12_1;
  assign _00595_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01959_ : lut_lookup_le_fraction_lpi_1_dfm_16_34_12_1;
  assign _00301_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) cfg_precision_1_sva_st_71 : cfg_precision_1_sva_st_107;
  assign _00445_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01970_ : lut_lookup_4_and_svs_2;
  assign _00645_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_lo_uflow_lpi_1_dfm_3 : lut_lookup_lo_uflow_lpi_1_dfm_4;
  assign _00419_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01969_ : lut_lookup_3_and_svs_2;
  assign _00643_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_lo_uflow_3_lpi_1_dfm_3 : lut_lookup_lo_uflow_3_lpi_1_dfm_4;
  assign _00394_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01968_ : lut_lookup_2_and_svs_2;
  assign _00641_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_lo_uflow_2_lpi_1_dfm_3 : lut_lookup_lo_uflow_2_lpi_1_dfm_4;
  assign _00369_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01967_ : lut_lookup_1_and_svs_2;
  assign _00639_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_lo_uflow_1_lpi_1_dfm_3 : lut_lookup_lo_uflow_1_lpi_1_dfm_4;
  assign _00646_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_else_unequal_tmp_18 : lut_lookup_unequal_tmp_13;
  assign _00357_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_in_data_sva_157 : lut_in_data_sva_158;
  assign _00266_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) cfg_lut_hybrid_priority_1_sva_9 : cfg_lut_hybrid_priority_1_sva_10;
  assign _00290_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) cfg_lut_oflow_priority_1_sva_9 : cfg_lut_oflow_priority_1_sva_10;
  assign _00295_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) cfg_lut_uflow_priority_1_sva_9 : cfg_lut_uflow_priority_1_sva_10;
  assign _00271_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) cfg_lut_le_function_1_sva_st_42 : cfg_lut_le_function_1_sva_10;
  assign _00602_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01979_ : lut_lookup_le_index_0_5_0_1_lpi_1_dfm_29;
  assign _00588_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01932_ : lut_lookup_le_fraction_1_lpi_1_dfm_22;
  assign _00601_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_le_index_0_5_0_1_lpi_1_dfm_27 : lut_lookup_le_index_0_5_0_1_lpi_1_dfm_28;
  assign _00587_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01934_ : lut_lookup_le_fraction_1_lpi_1_dfm_21;
  assign _00599_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_le_index_0_5_0_1_lpi_1_dfm_25 : lut_lookup_le_index_0_5_0_1_lpi_1_dfm_26;
  assign _00622_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01936_ : lut_lookup_lo_fraction_1_lpi_1_dfm_9;
  assign _00607_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01982_ : lut_lookup_le_index_0_5_0_2_lpi_1_dfm_29;
  assign _00591_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01942_ : lut_lookup_le_fraction_2_lpi_1_dfm_22;
  assign _00606_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_le_index_0_5_0_2_lpi_1_dfm_27 : lut_lookup_le_index_0_5_0_2_lpi_1_dfm_28;
  assign _00590_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01944_ : lut_lookup_le_fraction_2_lpi_1_dfm_21;
  assign _00604_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_le_index_0_5_0_2_lpi_1_dfm_25 : lut_lookup_le_index_0_5_0_2_lpi_1_dfm_26;
  assign _00623_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01946_ : lut_lookup_lo_fraction_2_lpi_1_dfm_9;
  assign _00612_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01976_ : lut_lookup_le_index_0_5_0_3_lpi_1_dfm_29;
  assign _00594_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01952_ : lut_lookup_le_fraction_3_lpi_1_dfm_22;
  assign _00611_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_le_index_0_5_0_3_lpi_1_dfm_27 : lut_lookup_le_index_0_5_0_3_lpi_1_dfm_28;
  assign _00593_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01954_ : lut_lookup_le_fraction_3_lpi_1_dfm_21;
  assign _00609_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_le_index_0_5_0_3_lpi_1_dfm_25 : lut_lookup_le_index_0_5_0_3_lpi_1_dfm_26;
  assign _00624_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01956_ : lut_lookup_lo_fraction_3_lpi_1_dfm_9;
  assign _00617_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01973_ : lut_lookup_le_index_0_5_0_lpi_1_dfm_29;
  assign _00597_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01962_ : lut_lookup_le_fraction_lpi_1_dfm_22;
  assign _00616_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_le_index_0_5_0_lpi_1_dfm_27 : lut_lookup_le_index_0_5_0_lpi_1_dfm_28;
  assign _00596_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01964_ : lut_lookup_le_fraction_lpi_1_dfm_21;
  assign _00614_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_le_index_0_5_0_lpi_1_dfm_25 : lut_lookup_le_index_0_5_0_lpi_1_dfm_26;
  assign _00625_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) _01966_ : lut_lookup_lo_fraction_lpi_1_dfm_9;
  assign _00544_ = cfg_lut_hybrid_priority_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9485" *) lut_lookup_else_unequal_tmp_12 : lut_lookup_else_unequal_tmp_13;
  assign _00651_ = _01926_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9433" *) _02590_ : main_stage_v_5;
  assign _00449_ = _01924_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9424" *) FpAdd_8U_23U_2_mux_61_itm_3 : lut_lookup_4_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  assign _00168_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9414" *) _02586_ : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_4_itm_1_0_1;
  assign _00437_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9414" *) nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 : lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  assign _00833_ = and_430_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_4_if_else_else_else_if_acc_nl[3] : FpAdd_8U_23U_1_mux_61_itm_4;
  assign _00502_ = _01923_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9404" *) _00833_ : lut_lookup_else_else_else_asn_mdf_sva_st_3;
  assign _00176_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9394" *) _02585_ : FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_4_itm_1_0_1;
  assign _00439_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9394" *) z_out_7[7:0] : lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  assign _00581_ = _01922_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9385" *) IsNaN_8U_23U_1_land_lpi_1_dfm_8 : lut_lookup_if_else_else_slc_10_mdf_sva_st_3;
  assign _00832_ = and_428_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_if_lor_1_lpi_1_dfm_mx0w1 : lut_lookup_4_if_else_else_else_else_acc_nl[32];
  assign _00452_ = _01921_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9375" *) _00832_ : lut_lookup_4_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _00423_ = _01920_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9364" *) FpAdd_8U_23U_2_mux_45_itm_3 : lut_lookup_3_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  assign _00167_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9354" *) _02586_ : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_3_itm_1_0_1;
  assign _00411_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9354" *) nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 : lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  assign _00831_ = and_430_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_3_if_else_else_else_if_acc_nl[3] : FpAdd_8U_23U_1_mux_45_itm_4;
  assign _00499_ = _01919_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9344" *) _00831_ : lut_lookup_else_else_else_asn_mdf_3_sva_st_3;
  assign _00175_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9334" *) _02585_ : FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_3_itm_1_0_1;
  assign _00413_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9334" *) z_out_6[7:0] : lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  assign _00578_ = _01918_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9325" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_8 : lut_lookup_if_else_else_slc_10_mdf_3_sva_st_3;
  assign _00830_ = and_428_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_if_lor_7_lpi_1_dfm_mx0w1 : lut_lookup_3_if_else_else_else_else_acc_nl[32];
  assign _00426_ = _01917_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9315" *) _00830_ : lut_lookup_3_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _00398_ = _01916_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9304" *) FpAdd_8U_23U_2_mux_29_itm_3 : lut_lookup_2_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  assign _00166_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9294" *) _02586_ : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_2_itm_1_0_1;
  assign _00386_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9294" *) nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 : lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  assign _00829_ = and_430_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_2_if_else_else_else_if_acc_nl[3] : FpAdd_8U_23U_1_mux_29_itm_4;
  assign _00496_ = _01915_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9284" *) _00829_ : lut_lookup_else_else_else_asn_mdf_2_sva_st_3;
  assign _00174_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9274" *) _02585_ : FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_2_itm_1_0_1;
  assign _00388_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9274" *) z_out_5[7:0] : lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  assign _00575_ = _01914_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9265" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_8 : lut_lookup_if_else_else_slc_10_mdf_2_sva_st_3;
  assign _00828_ = and_428_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_if_lor_6_lpi_1_dfm_mx0w1 : lut_lookup_2_if_else_else_else_else_acc_nl[32];
  assign _00401_ = _01913_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9255" *) _00828_ : lut_lookup_2_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _00373_ = _01912_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9244" *) FpAdd_8U_23U_2_mux_13_itm_3 : lut_lookup_1_else_1_else_if_slc_lut_lookup_else_1_else_lo_index_s_8_2_itm_3;
  assign _00169_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9234" *) _02586_ : FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_itm_1_0_1;
  assign _00361_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9234" *) nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2 : lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_abs_expo_acc_itm_2;
  assign _00827_ = and_430_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_1_if_else_else_else_if_acc_nl[3] : FpAdd_8U_23U_1_mux_13_itm_4;
  assign _00493_ = _01911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9224" *) _00827_ : lut_lookup_else_else_else_asn_mdf_1_sva_st_3;
  assign _00177_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9214" *) _02585_ : FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_1_0_1;
  assign _00363_ = FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9214" *) z_out_4[7:0] : lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_abs_expo_acc_itm_2;
  assign _00861_ = lut_lookup_else_else_slc_32_mdf_1_sva_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_1_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 : 6'b000000;
  assign _00860_ = lut_lookup_else_else_slc_32_mdf_2_sva_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_2_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 : 6'b000000;
  assign _00859_ = lut_lookup_else_else_slc_32_mdf_3_sva_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_3_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 : 6'b000000;
  assign _00858_ = lut_lookup_else_else_slc_32_mdf_sva_7 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13595|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13594" *) lut_lookup_4_if_else_else_else_else_slc_lut_lookup_if_else_else_else_le_index_s_5_0_itm_2 : 6'b000000;
  assign _00273_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) cfg_lut_le_function_1_sva_st_41 : cfg_lut_le_function_1_sva_st_42;
  assign _00303_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) cfg_precision_1_sva_st_70 : cfg_precision_1_sva_st_71;
  assign _00356_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) lut_in_data_sva_156 : lut_in_data_sva_157;
  assign _00270_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) cfg_lut_hybrid_priority_1_sva_8 : cfg_lut_hybrid_priority_1_sva_9;
  assign _00294_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) cfg_lut_oflow_priority_1_sva_8 : cfg_lut_oflow_priority_1_sva_9;
  assign _00299_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) cfg_lut_uflow_priority_1_sva_8 : cfg_lut_uflow_priority_1_sva_9;
  assign _00600_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) _01909_ : lut_lookup_le_index_0_5_0_1_lpi_1_dfm_27;
  assign _00598_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) _00861_ : lut_lookup_le_index_0_5_0_1_lpi_1_dfm_25;
  assign _00605_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) _01906_ : lut_lookup_le_index_0_5_0_2_lpi_1_dfm_27;
  assign _00603_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) _00860_ : lut_lookup_le_index_0_5_0_2_lpi_1_dfm_25;
  assign _00610_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) _01903_ : lut_lookup_le_index_0_5_0_3_lpi_1_dfm_27;
  assign _00608_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) _00859_ : lut_lookup_le_index_0_5_0_3_lpi_1_dfm_25;
  assign _00615_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) _01900_ : lut_lookup_le_index_0_5_0_lpi_1_dfm_27;
  assign _00613_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) _00858_ : lut_lookup_le_index_0_5_0_lpi_1_dfm_25;
  assign _00545_ = cfg_precision_and_24_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9175" *) lut_lookup_unequal_tmp_mx0w0 : lut_lookup_else_unequal_tmp_18;
  assign _00458_ = lut_lookup_if_else_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9150" *) FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6 : lut_lookup_4_if_else_slc_32_svs_st_5;
  assign _00432_ = lut_lookup_if_else_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9150" *) FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6 : lut_lookup_3_if_else_slc_32_svs_st_5;
  assign _00407_ = lut_lookup_if_else_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9150" *) FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6 : lut_lookup_2_if_else_slc_32_svs_st_5;
  assign _00382_ = lut_lookup_if_else_if_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9150" *) FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6 : lut_lookup_1_if_else_slc_32_svs_st_5;
  assign _00572_ = _01897_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9139" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_8 : lut_lookup_if_else_else_slc_10_mdf_1_sva_st_3;
  assign _00826_ = and_428_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_if_lor_5_lpi_1_dfm_mx0w1 : lut_lookup_1_if_else_else_else_else_acc_nl[32];
  assign _00376_ = _01896_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9129" *) _00826_ : lut_lookup_1_if_else_else_else_else_if_slc_lut_lookup_if_else_else_else_else_acc_32_svs_st_2;
  assign _00277_ = _00924_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9119" *) cfg_lut_le_index_offset_1_sva_6 : cfg_lut_le_index_offset_1_sva_7;
  assign _00650_ = _01895_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9111" *) _02580_ : main_stage_v_4;
  assign _00825_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : FpAdd_8U_23U_2_mux_61_itm_1;
  assign _00149_ = _01893_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9102" *) _00825_ : FpAdd_8U_23U_2_mux_61_itm_3;
  assign _00153_ = _01892_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9090" *) _03314_ : FpAdd_8U_23U_2_o_expo_lpi_1_dfm_12;
  assign _00824_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : FpMantRNE_49U_24U_2_else_carry_sva_mx0w0;
  assign _00189_ = _01890_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9078" *) _00824_ : FpMantRNE_49U_24U_2_else_carry_sva_2;
  assign _00443_ = _01889_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9068" *) FpAdd_8U_23U_2_int_mant_1_lpi_1_dfm_2_mx0[47:25] : lut_lookup_4_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  assign _00823_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_4_else_else_else_if_acc_nl[3] : FpAdd_8U_23U_1_mux_61_itm_3;
  assign _00117_ = _01888_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9057" *) _00823_ : FpAdd_8U_23U_1_mux_61_itm_4;
  assign _00658_ = _01887_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9047" *) _03286_ : reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm;
  assign _00659_ = _01885_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9037" *) _03266_ : reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_itm;
  assign _00441_ = FpMantRNE_49U_24U_1_else_o_mant_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9025" *) FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[47:25] : lut_lookup_4_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  assign _00185_ = FpMantRNE_49U_24U_1_else_o_mant_and_3_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9025" *) FpMantRNE_49U_24U_1_else_carry_sva_mx0w0 : FpMantRNE_49U_24U_1_else_carry_sva_2;
  assign _00725_ = _01882_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9014" *) lut_lookup_if_else_else_else_le_index_s_sva[7:6] : reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  assign _00726_ = _01878_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:9003" *) lut_lookup_if_else_else_else_le_index_s_sva[8] : reg_lut_lookup_4_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  assign _00212_ = _01877_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8992" *) _03192_ : IsNaN_8U_23U_1_land_lpi_1_dfm_8;
  assign _00822_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : FpAdd_8U_23U_2_mux_45_itm_1;
  assign _00146_ = _01876_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8982" *) _00822_ : FpAdd_8U_23U_2_mux_45_itm_3;
  assign _00152_ = _01875_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8970" *) _03313_ : FpAdd_8U_23U_2_o_expo_3_lpi_1_dfm_12;
  assign _00821_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : FpMantRNE_49U_24U_2_else_carry_3_sva_mx0w0;
  assign _00188_ = _01873_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8958" *) _00821_ : FpMantRNE_49U_24U_2_else_carry_3_sva_2;
  assign _00417_ = _01872_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8948" *) FpAdd_8U_23U_2_int_mant_4_lpi_1_dfm_2_mx0[47:25] : lut_lookup_3_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  assign _00820_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_3_else_else_else_if_acc_nl[3] : FpAdd_8U_23U_1_mux_45_itm_3;
  assign _00114_ = _01871_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8937" *) _00820_ : FpAdd_8U_23U_1_mux_45_itm_4;
  assign _00656_ = _01870_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8927" *) _03285_ : reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm;
  assign _00657_ = _01868_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8917" *) _03265_ : reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_itm;
  assign _00415_ = FpMantRNE_49U_24U_1_else_o_mant_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8905" *) FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[47:25] : lut_lookup_3_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  assign _00184_ = FpMantRNE_49U_24U_1_else_o_mant_and_2_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8905" *) FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w0 : FpMantRNE_49U_24U_1_else_carry_3_sva_2;
  assign _00714_ = _01865_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8894" *) lut_lookup_if_else_else_else_le_index_s_3_sva[7:6] : reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  assign _00715_ = _01861_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8883" *) lut_lookup_if_else_else_else_le_index_s_3_sva[8] : reg_lut_lookup_3_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  assign _00209_ = _01860_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8872" *) _03191_ : IsNaN_8U_23U_1_land_3_lpi_1_dfm_8;
  assign _00819_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : FpAdd_8U_23U_2_mux_29_itm_1;
  assign _00143_ = _01859_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8862" *) _00819_ : FpAdd_8U_23U_2_mux_29_itm_3;
  assign _00246_ = IsNaN_8U_23U_8_aelse_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8850" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5 : IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_6;
  assign _00244_ = IsNaN_8U_23U_8_aelse_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8850" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 : IsNaN_8U_23U_7_land_2_lpi_1_dfm_7;
  assign _00391_ = IsNaN_8U_23U_8_aelse_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8850" *) lut_lookup_2_FpMantRNE_49U_24U_2_else_and_tmp : lut_lookup_2_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign _00259_ = IsNaN_8U_23U_8_aelse_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8850" *) IsNaN_8U_23U_8_land_1_lpi_1_dfm_6 : IsNaN_8U_23U_8_land_2_lpi_1_dfm_7;
  assign _00151_ = _01858_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8836" *) _03312_ : FpAdd_8U_23U_2_o_expo_2_lpi_1_dfm_12;
  assign _00818_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : FpMantRNE_49U_24U_2_else_carry_2_sva_mx0w0;
  assign _00187_ = _01856_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8824" *) _00818_ : FpMantRNE_49U_24U_2_else_carry_2_sva_2;
  assign _00392_ = _01855_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8814" *) FpAdd_8U_23U_2_int_mant_3_lpi_1_dfm_2_mx0[47:25] : lut_lookup_2_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  assign _00817_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_1_land_lpi_1_dfm_7 : nor_50_cse_1;
  assign _00816_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_1_land_3_lpi_1_dfm_7 : nor_38_cse_1;
  assign _00815_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_7 : nor_27_cse_1;
  assign _00105_ = FpAdd_8U_23U_2_is_inf_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8800" *) _00817_ : FpAdd_8U_23U_1_is_inf_lpi_1_dfm_6;
  assign _00104_ = FpAdd_8U_23U_2_is_inf_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8800" *) _00816_ : FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_6;
  assign _00103_ = FpAdd_8U_23U_2_is_inf_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8800" *) _00815_ : FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_6;
  assign _00814_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_2_else_else_else_if_acc_nl[3] : FpAdd_8U_23U_1_mux_29_itm_3;
  assign _00111_ = _01854_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8788" *) _00814_ : FpAdd_8U_23U_1_mux_29_itm_4;
  assign _00654_ = _01853_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8778" *) _03284_ : reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm;
  assign _00655_ = _01851_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8768" *) _03264_ : reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_itm;
  assign _00390_ = FpMantRNE_49U_24U_1_else_o_mant_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8757" *) FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[47:25] : lut_lookup_2_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  assign _00183_ = FpMantRNE_49U_24U_1_else_o_mant_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8757" *) FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w0 : FpMantRNE_49U_24U_1_else_carry_2_sva_2;
  assign _00703_ = _01848_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8746" *) lut_lookup_if_else_else_else_le_index_s_2_sva[7:6] : reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  assign _00704_ = _01844_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8735" *) lut_lookup_if_else_else_else_le_index_s_2_sva[8] : reg_lut_lookup_2_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  assign _00207_ = _01843_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8724" *) _03190_ : IsNaN_8U_23U_1_land_2_lpi_1_dfm_8;
  assign _00813_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_7_land_lpi_1_dfm_6 : nor_54_cse;
  assign _00812_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 : nor_42_cse;
  assign _00811_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_6 : nor_31_cse;
  assign _00810_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 : nor_13_cse;
  assign _00137_ = FpAdd_8U_23U_2_is_inf_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8708" *) _00813_ : FpAdd_8U_23U_2_is_inf_lpi_1_dfm_5;
  assign _00136_ = FpAdd_8U_23U_2_is_inf_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8708" *) _00812_ : FpAdd_8U_23U_2_is_inf_3_lpi_1_dfm_5;
  assign _00135_ = FpAdd_8U_23U_2_is_inf_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8708" *) _00811_ : FpAdd_8U_23U_2_is_inf_2_lpi_1_dfm_5;
  assign _00134_ = FpAdd_8U_23U_2_is_inf_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8708" *) _00810_ : FpAdd_8U_23U_2_is_inf_1_lpi_1_dfm_5;
  assign _00809_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : FpAdd_8U_23U_2_mux_13_itm_1;
  assign _00139_ = _01841_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8696" *) _00809_ : FpAdd_8U_23U_2_mux_13_itm_3;
  assign _00288_ = _01840_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8687" *) cfg_lut_lo_start_1_sva_2_30_0_1 : cfg_lut_lo_start_1_sva_3_30_0_1;
  assign _00150_ = _01839_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8676" *) _03311_ : FpAdd_8U_23U_2_o_expo_1_lpi_1_dfm_12;
  assign _00808_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_obits_fixed_or_tmp[8] : FpMantRNE_49U_24U_2_else_carry_1_sva_mx0w0;
  assign _00186_ = _01837_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8665" *) _00808_ : FpMantRNE_49U_24U_2_else_carry_1_sva_2;
  assign _00367_ = _01836_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8655" *) FpAdd_8U_23U_2_int_mant_2_lpi_1_dfm_2_mx0[47:25] : lut_lookup_1_FpMantRNE_49U_24U_2_else_o_mant_slc_FpMantRNE_49U_24U_i_data_2_48_25_2_itm_2;
  assign _00807_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_1_land_1_lpi_1_dfm_7 : nor_5_cse_1;
  assign _00102_ = _01835_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8645" *) _00807_ : FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_6;
  assign _00718_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) lut_lookup_4_FpMantRNE_49U_24U_else_and_tmp : reg_lut_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign _00707_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) lut_lookup_3_FpMantRNE_49U_24U_else_and_tmp : reg_lut_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign _00696_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) lut_lookup_2_FpMantRNE_49U_24U_else_and_tmp : reg_lut_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign _00685_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) lut_lookup_1_FpMantRNE_49U_24U_else_and_tmp : reg_lut_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign _00254_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse : IsNaN_8U_23U_7_land_lpi_1_dfm_st_6;
  assign _00251_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5 : IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_6;
  assign _00242_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5 : IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_6;
  assign _00253_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) IsNaN_8U_23U_7_land_lpi_1_dfm_6 : IsNaN_8U_23U_7_land_lpi_1_dfm_7;
  assign _00442_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) lut_lookup_4_FpMantRNE_49U_24U_2_else_and_tmp : lut_lookup_4_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign _00248_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_6 : IsNaN_8U_23U_7_land_3_lpi_1_dfm_7;
  assign _00416_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) lut_lookup_3_FpMantRNE_49U_24U_2_else_and_tmp : lut_lookup_3_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign _00239_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_6 : IsNaN_8U_23U_7_land_1_lpi_1_dfm_7;
  assign _00366_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) lut_lookup_1_FpMantRNE_49U_24U_2_else_and_tmp : lut_lookup_1_FpMantRNE_49U_24U_2_else_and_svs_2;
  assign _00261_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) IsNaN_8U_23U_8_land_3_lpi_1_dfm_4 : IsNaN_8U_23U_8_land_3_lpi_1_dfm_5;
  assign _00263_ = FpMantRNE_49U_24U_1_else_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8622" *) IsNaN_8U_23U_8_land_lpi_1_dfm_4 : IsNaN_8U_23U_8_land_lpi_1_dfm_5;
  assign _00806_ = and_dcpl_162 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_4_land_lpi_1_dfm_4 : reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse;
  assign _00805_ = and_dcpl_162 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse : IsNaN_8U_23U_1_land_lpi_1_dfm_7;
  assign _00804_ = and_dcpl_162 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_4_land_3_lpi_1_dfm_5 : IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5;
  assign _00803_ = and_dcpl_162 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5 : IsNaN_8U_23U_1_land_3_lpi_1_dfm_7;
  assign _00802_ = and_dcpl_162 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_4_land_2_lpi_1_dfm_5 : IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5;
  assign _00801_ = and_dcpl_162 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5 : IsNaN_8U_23U_1_land_2_lpi_1_dfm_7;
  assign _00800_ = and_dcpl_162 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_4_land_1_lpi_1_dfm_4 : IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5;
  assign _00799_ = and_dcpl_162 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5 : IsNaN_8U_23U_1_land_1_lpi_1_dfm_7;
  assign _00221_ = IsNaN_8U_23U_3_aelse_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8584" *) _00806_ : IsNaN_8U_23U_3_land_lpi_1_dfm_st_6;
  assign _00219_ = IsNaN_8U_23U_3_aelse_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8584" *) _00804_ : IsNaN_8U_23U_3_land_3_lpi_1_dfm_st_6;
  assign _00217_ = IsNaN_8U_23U_3_aelse_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8584" *) _00802_ : IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_6;
  assign _00214_ = IsNaN_8U_23U_3_aelse_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8584" *) _00800_ : IsNaN_8U_23U_3_land_1_lpi_1_dfm_st_6;
  assign _00220_ = IsNaN_8U_23U_3_aelse_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8584" *) _00805_ : IsNaN_8U_23U_3_land_lpi_1_dfm_6;
  assign _00218_ = IsNaN_8U_23U_3_aelse_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8584" *) _00803_ : IsNaN_8U_23U_3_land_3_lpi_1_dfm_7;
  assign _00215_ = IsNaN_8U_23U_3_aelse_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8584" *) _00801_ : IsNaN_8U_23U_3_land_2_lpi_1_dfm_7;
  assign _00213_ = IsNaN_8U_23U_3_aelse_and_6_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8584" *) _00799_ : IsNaN_8U_23U_3_land_1_lpi_1_dfm_6;
  assign _00798_ = and_dcpl_161 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_1_else_else_else_if_acc_nl[3] : FpAdd_8U_23U_1_mux_13_itm_3;
  assign _00107_ = _01834_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8568" *) _00798_ : FpAdd_8U_23U_1_mux_13_itm_4;
  assign _00652_ = _01832_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8558" *) _03283_ : reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm;
  assign _00653_ = _01830_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8548" *) _03263_ : reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_itm;
  assign _00365_ = FpMantRNE_49U_24U_1_else_o_mant_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8537" *) FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[47:25] : lut_lookup_1_FpMantRNE_49U_24U_1_else_o_mant_slc_FpMantRNE_49U_24U_i_data_1_48_25_2_itm_2;
  assign _00182_ = FpMantRNE_49U_24U_1_else_o_mant_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8537" *) FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w0 : FpMantRNE_49U_24U_1_else_carry_1_sva_2;
  assign _00692_ = _01827_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8526" *) lut_lookup_if_else_else_else_le_index_s_1_sva[7:6] : reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_1_itm;
  assign _00693_ = _01823_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8515" *) lut_lookup_if_else_else_else_le_index_s_1_sva[8] : reg_lut_lookup_1_if_else_else_else_if_slc_lut_lookup_if_else_else_else_le_index_s_8_6_itm;
  assign _00204_ = _01822_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8504" *) _03189_ : IsNaN_8U_23U_1_land_1_lpi_1_dfm_8;
  assign _00282_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) cfg_lut_le_start_1_sva_2_30_0_1 : cfg_lut_le_start_1_sva_3_30_0_1;
  assign _00272_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) reg_cfg_lut_le_function_1_sva_st_20_cse : cfg_lut_le_function_1_sva_st_41;
  assign _00302_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) reg_cfg_precision_1_sva_st_13_cse_1 : cfg_precision_1_sva_st_70;
  assign _00355_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) lut_in_data_sva_155 : lut_in_data_sva_156;
  assign _00269_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) cfg_lut_hybrid_priority_1_sva_7 : cfg_lut_hybrid_priority_1_sva_8;
  assign _00293_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) cfg_lut_oflow_priority_1_sva_7 : cfg_lut_oflow_priority_1_sva_8;
  assign _00298_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) cfg_lut_uflow_priority_1_sva_7 : cfg_lut_uflow_priority_1_sva_8;
  assign _00286_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) cfg_lut_lo_index_select_1_sva_5 : cfg_lut_lo_index_select_1_sva_6;
  assign _00280_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) cfg_lut_le_index_select_1_sva_5 : cfg_lut_le_index_select_1_sva_6;
  assign _00276_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) cfg_lut_le_index_offset_1_sva_5 : cfg_lut_le_index_offset_1_sva_6;
  assign _00570_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) lut_lookup_1_if_else_else_acc_nl[10] : lut_lookup_if_else_else_slc_10_mdf_1_sva_3;
  assign _00573_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) lut_lookup_2_if_else_else_acc_nl[10] : lut_lookup_if_else_else_slc_10_mdf_2_sva_3;
  assign _00576_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) lut_lookup_3_if_else_else_acc_nl[10] : lut_lookup_if_else_else_slc_10_mdf_3_sva_3;
  assign _00579_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) lut_lookup_4_if_else_else_acc_nl[10] : lut_lookup_if_else_else_slc_10_mdf_sva_3;
  assign _00380_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) lut_lookup_1_if_else_slc_32_svs_6 : lut_lookup_1_if_else_slc_32_svs_7;
  assign _00405_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) lut_lookup_2_if_else_slc_32_svs_6 : lut_lookup_2_if_else_slc_32_svs_7;
  assign _00430_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) lut_lookup_3_if_else_slc_32_svs_6 : lut_lookup_3_if_else_slc_32_svs_7;
  assign _00456_ = cfg_lut_le_start_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8478" *) lut_lookup_4_if_else_slc_32_svs_6 : lut_lookup_4_if_else_slc_32_svs_7;
  assign _00649_ = _01820_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8453" *) _02556_ : main_stage_v_3;
  assign _00853_ = and_338_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13578|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13577" *) lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl : lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl;
  assign _00129_ = _01818_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8444" *) _00853_ : FpAdd_8U_23U_2_int_mant_p1_sva_3;
  assign _00097_ = _01815_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8432" *) _03278_ : FpAdd_8U_23U_1_int_mant_p1_sva_3;
  assign _00666_ = _01813_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8423" *) FpAdd_8U_23U_1_mux1h_7_itm[5:0] : reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm;
  assign _00852_ = and_324_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13578|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13577" *) lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl : lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl;
  assign _00128_ = _01810_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8413" *) _00852_ : FpAdd_8U_23U_2_int_mant_p1_3_sva_3;
  assign _00677_ = FpAdd_8U_23U_2_and_37_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8399" *) reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse : reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_2_cse;
  assign _00250_ = FpAdd_8U_23U_2_and_37_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8399" *) IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4 : IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_5;
  assign _00165_ = FpAdd_8U_23U_2_and_37_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8399" *) FpAdd_8U_23U_2_qr_lpi_1_dfm_4 : FpAdd_8U_23U_2_qr_lpi_1_dfm_5;
  assign _00163_ = FpAdd_8U_23U_2_and_37_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8399" *) FpAdd_8U_23U_2_qr_4_lpi_1_dfm_4 : FpAdd_8U_23U_2_qr_4_lpi_1_dfm_5;
  assign _00260_ = FpAdd_8U_23U_2_and_37_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8399" *) nor_482_cse : IsNaN_8U_23U_8_land_3_lpi_1_dfm_4;
  assign _00262_ = FpAdd_8U_23U_2_and_37_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8399" *) nor_469_cse : IsNaN_8U_23U_8_land_lpi_1_dfm_4;
  assign _00096_ = _01807_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8383" *) _03277_ : FpAdd_8U_23U_1_int_mant_p1_3_sva_3;
  assign _00664_ = _01805_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8374" *) FpAdd_8U_23U_1_mux1h_5_itm[5:0] : reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm;
  assign _00851_ = and_308_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13578|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13577" *) lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl : lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl;
  assign _00127_ = _01802_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8364" *) _00851_ : FpAdd_8U_23U_2_int_mant_p1_2_sva_3;
  assign _00245_ = FpAdd_8U_23U_2_and_36_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8354" *) IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4 : IsNaN_8U_23U_7_land_2_lpi_1_dfm_st_5;
  assign _00161_ = FpAdd_8U_23U_2_and_36_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8354" *) FpAdd_8U_23U_2_qr_3_lpi_1_dfm_4 : FpAdd_8U_23U_2_qr_3_lpi_1_dfm_5;
  assign _00095_ = _01799_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8342" *) _03276_ : FpAdd_8U_23U_1_int_mant_p1_2_sva_3;
  assign _00662_ = _01797_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8333" *) FpAdd_8U_23U_1_mux1h_3_itm[5:0] : reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm;
  assign _00667_ = and_961_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8322" *) FpAdd_8U_23U_1_mux1h_7_itm[7:6] : reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_itm;
  assign _00665_ = and_961_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8322" *) FpAdd_8U_23U_1_mux1h_5_itm[7:6] : reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_itm;
  assign _00663_ = and_961_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8322" *) FpAdd_8U_23U_1_mux1h_3_itm[7:6] : reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_itm;
  assign _00850_ = and_292_rgt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13578|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13577" *) lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl : lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl;
  assign _00126_ = _01794_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8311" *) _00850_ : FpAdd_8U_23U_2_int_mant_p1_1_sva_3;
  assign _00241_ = FpAdd_8U_23U_2_and_35_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8300" *) IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4 : IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_5;
  assign _00159_ = FpAdd_8U_23U_2_and_35_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8300" *) FpAdd_8U_23U_2_qr_2_lpi_1_dfm_4 : FpAdd_8U_23U_2_qr_2_lpi_1_dfm_5;
  assign _00257_ = FpAdd_8U_23U_2_and_35_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8300" *) IsNaN_8U_23U_8_land_2_lpi_1_dfm_5 : IsNaN_8U_23U_8_land_1_lpi_1_dfm_6;
  assign _00094_ = _01791_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8287" *) _03275_ : FpAdd_8U_23U_1_int_mant_p1_1_sva_3;
  assign _00660_ = _01789_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8278" *) FpAdd_8U_23U_1_mux1h_1_itm[5:0] : reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm;
  assign _00661_ = _01786_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8269" *) FpAdd_8U_23U_1_mux1h_1_itm[7:6] : reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_itm;
  assign _00679_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) reg_cfg_lut_le_function_1_sva_st_19_cse : reg_cfg_lut_le_function_1_sva_st_20_cse;
  assign _00681_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) reg_cfg_precision_1_sva_st_12_cse_1 : reg_cfg_precision_1_sva_st_13_cse_1;
  assign _00287_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) cfg_lut_lo_start_1_sva_41[30:0] : cfg_lut_lo_start_1_sva_2_30_0_1;
  assign _00281_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) cfg_lut_le_start_1_sva_41[30:0] : cfg_lut_le_start_1_sva_2_30_0_1;
  assign _00354_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) lut_in_data_sva_154 : lut_in_data_sva_155;
  assign _00268_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) cfg_lut_hybrid_priority_1_sva_6 : cfg_lut_hybrid_priority_1_sva_7;
  assign _00292_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) cfg_lut_oflow_priority_1_sva_6 : cfg_lut_oflow_priority_1_sva_7;
  assign _00297_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) cfg_lut_uflow_priority_1_sva_6 : cfg_lut_uflow_priority_1_sva_7;
  assign _00285_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) cfg_lut_lo_index_select_1_sva_4 : cfg_lut_lo_index_select_1_sva_5;
  assign _00279_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) cfg_lut_le_index_select_1_sva_4 : cfg_lut_le_index_select_1_sva_5;
  assign _00275_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) cfg_lut_le_index_offset_1_sva_4 : cfg_lut_le_index_offset_1_sva_5;
  assign _00379_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) lut_lookup_1_if_else_slc_32_svs_5 : lut_lookup_1_if_else_slc_32_svs_6;
  assign _00404_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) lut_lookup_2_if_else_slc_32_svs_5 : lut_lookup_2_if_else_slc_32_svs_6;
  assign _00429_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) lut_lookup_3_if_else_slc_32_svs_5 : lut_lookup_3_if_else_slc_32_svs_6;
  assign _00455_ = cfg_lut_le_index_offset_and_1_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8246" *) lut_lookup_4_if_else_slc_32_svs_5 : lut_lookup_4_if_else_slc_32_svs_6;
  assign _00648_ = _01783_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8224" *) _02551_ : main_stage_v_2;
  assign _00869_ = and_dcpl_304 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) cfg_lut_le_start_rsci_d[30:23] : chn_lut_in_rsci_d_mxwt[126:119];
  assign _00868_ = and_dcpl_296 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) cfg_lut_le_start_rsci_d[30:23] : chn_lut_in_rsci_d_mxwt[94:87];
  assign _00867_ = and_dcpl_288 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) cfg_lut_le_start_rsci_d[30:23] : chn_lut_in_rsci_d_mxwt[62:55];
  assign _00676_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0 : reg_IsNaN_8U_23U_3_land_lpi_1_dfm_st_1_cse;
  assign _00717_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _03913_ : reg_lut_lookup_4_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign _00716_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _03912_ : reg_lut_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign _00706_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _03911_ : reg_lut_lookup_3_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign _00705_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _03910_ : reg_lut_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign _00694_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _03908_ : reg_lut_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign _00695_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _03909_ : reg_lut_lookup_2_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign _00249_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _02548_ : IsNaN_8U_23U_7_land_3_lpi_1_dfm_st_4;
  assign _00216_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _02549_ : IsNaN_8U_23U_3_land_2_lpi_1_dfm_st_4;
  assign _00385_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) lut_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 : lut_lookup_2_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  assign _00121_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _00869_ : FpAdd_8U_23U_1_qr_lpi_1_dfm_5;
  assign _00120_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _00868_ : FpAdd_8U_23U_1_qr_4_lpi_1_dfm_5;
  assign _00119_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _00867_ : FpAdd_8U_23U_1_qr_3_lpi_1_dfm_5;
  assign _00091_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) acc_8_nl[8:1] : FpAdd_8U_23U_1_a_right_shift_qr_2_sva_3;
  assign _00092_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) acc_11_nl[8:1] : FpAdd_8U_23U_1_a_right_shift_qr_3_sva_3;
  assign _00093_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) acc_7_nl[8:1] : FpAdd_8U_23U_1_a_right_shift_qr_sva_3;
  assign _00205_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) IsNaN_8U_23U_1_land_2_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_1_land_2_lpi_1_dfm_6;
  assign _00258_ = FpAdd_8U_23U_1_is_addition_and_1_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8190" *) _02550_ : IsNaN_8U_23U_8_land_2_lpi_1_dfm_5;
  assign _00866_ = and_dcpl_284 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13612|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13611" *) cfg_lut_lo_start_rsci_d[30:23] : chn_lut_in_rsci_d_mxwt[30:23];
  assign _00684_ = FpAdd_8U_23U_2_is_addition_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8153" *) _03907_ : reg_lut_lookup_1_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_FpAdd_8U_23U_2_is_addition_xor_svs_st_1_cse;
  assign _00240_ = FpAdd_8U_23U_2_is_addition_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8153" *) IsNaN_8U_23U_3_land_1_lpi_1_dfm_mx0w0 : IsNaN_8U_23U_7_land_1_lpi_1_dfm_st_4;
  assign _00360_ = FpAdd_8U_23U_2_is_addition_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8153" *) lut_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_mx0w1 : lut_lookup_1_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2;
  assign _00158_ = FpAdd_8U_23U_2_is_addition_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8153" *) _00866_ : FpAdd_8U_23U_2_qr_2_lpi_1_dfm_4;
  assign _00122_ = FpAdd_8U_23U_2_is_addition_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8153" *) acc_6_nl[8:1] : FpAdd_8U_23U_2_a_right_shift_qr_1_sva_3;
  assign _00683_ = _01781_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8139" *) _03906_ : reg_lut_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_1_cse;
  assign _00678_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) cfg_lut_le_function_rsci_d : reg_cfg_lut_le_function_1_sva_st_19_cse;
  assign _00680_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) cfg_precision_rsci_d : reg_cfg_precision_1_sva_st_12_cse_1;
  assign _00353_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) chn_lut_in_rsci_d_mxwt : lut_in_data_sva_154;
  assign _00267_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) cfg_lut_hybrid_priority_rsci_d : cfg_lut_hybrid_priority_1_sva_6;
  assign _00291_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) cfg_lut_oflow_priority_rsci_d : cfg_lut_oflow_priority_1_sva_6;
  assign _00296_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) cfg_lut_uflow_priority_rsci_d : cfg_lut_uflow_priority_1_sva_6;
  assign _00284_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) cfg_lut_lo_index_select_rsci_d : cfg_lut_lo_index_select_1_sva_4;
  assign _00278_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) cfg_lut_le_index_select_rsci_d : cfg_lut_le_index_select_1_sva_4;
  assign _00274_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) cfg_lut_le_index_offset_rsci_d : cfg_lut_le_index_offset_1_sva_4;
  assign _00289_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) cfg_lut_lo_start_rsci_d : cfg_lut_lo_start_1_sva_41;
  assign _00283_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) cfg_lut_le_start_rsci_d : cfg_lut_le_start_1_sva_41;
  assign _00378_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) lut_lookup_1_else_else_acc_1_nl[32] : lut_lookup_1_if_else_slc_32_svs_5;
  assign _00403_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) lut_lookup_2_else_else_acc_1_nl[32] : lut_lookup_2_if_else_slc_32_svs_5;
  assign _00428_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) lut_lookup_3_else_else_acc_1_nl[32] : lut_lookup_3_if_else_slc_32_svs_5;
  assign _00454_ = cfg_precision_and_cse ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8116" *) lut_lookup_4_else_else_acc_1_nl[32] : lut_lookup_4_if_else_slc_32_svs_5;
  assign _00647_ = _01780_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8094" *) _02547_ : main_stage_v_1;
  assign _00682_ = _01779_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8086" *) _02546_ : reg_chn_lut_out_rsci_ld_core_psct_cse;
  assign _00797_ = and_dcpl_71 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_118_nl : lut_lookup_if_2_lut_lookup_if_2_and_15_nl;
  assign _00796_ = and_dcpl_71 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_117_nl : lut_lookup_if_2_lut_lookup_if_2_and_14_nl;
  assign _00795_ = and_dcpl_71 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_116_nl : lut_lookup_if_2_mux_24_nl;
  assign _00794_ = and_dcpl_71 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_106_nl : cfg_lut_uflow_priority_1_sva_10;
  assign _00793_ = and_dcpl_71 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_lut_lookup_else_2_and_7_nl : lut_lookup_else_2_else_else_if_mux_26_itm_1;
  assign _00319_ = chn_lut_out_and_16_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8069" *) _00793_ : chn_lut_out_rsci_d_275;
  assign _00323_ = chn_lut_out_and_16_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8069" *) _00794_ : chn_lut_out_rsci_d_279;
  assign _00337_ = chn_lut_out_and_16_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8069" *) _00795_ : chn_lut_out_rsci_d_313;
  assign _00338_ = chn_lut_out_and_16_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8069" *) _00796_ : chn_lut_out_rsci_d_314;
  assign _00339_ = chn_lut_out_and_16_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8069" *) _00797_ : chn_lut_out_rsci_d_315;
  assign _00792_ = and_dcpl_67 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_115_nl : lut_lookup_if_2_lut_lookup_if_2_and_13_nl;
  assign _00791_ = and_dcpl_67 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_114_nl : lut_lookup_if_2_lut_lookup_if_2_and_12_nl;
  assign _00790_ = and_dcpl_67 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_113_nl : lut_lookup_if_2_mux_23_nl;
  assign _00789_ = and_dcpl_67 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_105_nl : cfg_lut_uflow_priority_1_sva_10;
  assign _00788_ = and_dcpl_67 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_lut_lookup_else_2_and_6_nl : lut_lookup_else_2_else_else_if_mux_19_itm_1;
  assign _00318_ = chn_lut_out_and_15_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8048" *) _00788_ : chn_lut_out_rsci_d_274;
  assign _00322_ = chn_lut_out_and_15_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8048" *) _00789_ : chn_lut_out_rsci_d_278;
  assign _00333_ = chn_lut_out_and_15_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8048" *) _00790_ : chn_lut_out_rsci_d_304;
  assign _00334_ = chn_lut_out_and_15_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8048" *) _00791_ : chn_lut_out_rsci_d_305;
  assign _00335_ = chn_lut_out_and_15_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8048" *) _00792_ : chn_lut_out_rsci_d_306;
  assign _00787_ = and_dcpl_63 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_112_nl : lut_lookup_if_2_lut_lookup_if_2_and_11_nl;
  assign _00786_ = and_dcpl_63 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_111_nl : lut_lookup_if_2_lut_lookup_if_2_and_10_nl;
  assign _00785_ = and_dcpl_63 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_110_nl : lut_lookup_if_2_mux_22_nl;
  assign _00784_ = and_dcpl_63 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_104_nl : cfg_lut_uflow_priority_1_sva_10;
  assign _00783_ = and_dcpl_63 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_lut_lookup_else_2_and_5_nl : lut_lookup_else_2_else_else_if_mux_12_itm_1;
  assign _00317_ = chn_lut_out_and_14_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8027" *) _00783_ : chn_lut_out_rsci_d_273;
  assign _00321_ = chn_lut_out_and_14_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8027" *) _00784_ : chn_lut_out_rsci_d_277;
  assign _00329_ = chn_lut_out_and_14_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8027" *) _00785_ : chn_lut_out_rsci_d_295;
  assign _00330_ = chn_lut_out_and_14_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8027" *) _00786_ : chn_lut_out_rsci_d_296;
  assign _00331_ = chn_lut_out_and_14_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8027" *) _00787_ : chn_lut_out_rsci_d_297;
  assign _00782_ = and_dcpl_59 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_109_nl : lut_lookup_if_2_lut_lookup_if_2_and_9_nl;
  assign _00781_ = and_dcpl_59 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_108_nl : lut_lookup_if_2_lut_lookup_if_2_and_8_nl;
  assign _00780_ = and_dcpl_59 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_107_nl : lut_lookup_if_2_mux_21_nl;
  assign _00779_ = and_dcpl_59 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_mux_103_nl : cfg_lut_uflow_priority_1_sva_10;
  assign _00778_ = and_dcpl_59 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13459|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13458" *) lut_lookup_else_2_lut_lookup_else_2_and_4_nl : lut_lookup_else_2_else_else_if_mux_5_itm_1;
  assign _00316_ = chn_lut_out_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8006" *) _00778_ : chn_lut_out_rsci_d_272;
  assign _00320_ = chn_lut_out_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8006" *) _00779_ : chn_lut_out_rsci_d_276;
  assign _00325_ = chn_lut_out_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8006" *) _00780_ : chn_lut_out_rsci_d_286;
  assign _00326_ = chn_lut_out_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8006" *) _00781_ : chn_lut_out_rsci_d_287;
  assign _00327_ = chn_lut_out_and_13_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8006" *) _00782_ : chn_lut_out_rsci_d_288;
  assign _00845_ = lut_lookup_not_36_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13476|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13475" *) lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_4_nl : 12'b000000000000;
  assign _00844_ = lut_lookup_not_37_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13476|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13475" *) lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_5_nl : 12'b000000000000;
  assign _00843_ = lut_lookup_not_38_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13476|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13475" *) lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_6_nl : 12'b000000000000;
  assign _00842_ = lut_lookup_not_39_nl ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13476|./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:13475" *) lut_lookup_lut_lookup_lut_lookup_lut_lookup_mux1h_7_nl : 12'b000000000000;
  assign _00309_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _00842_ : chn_lut_out_rsci_d_11_0;
  assign _00348_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _03255_ : chn_lut_out_rsci_d_34_12;
  assign _00349_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _00843_ : chn_lut_out_rsci_d_46_35;
  assign _00350_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _03256_ : chn_lut_out_rsci_d_69_47;
  assign _00351_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _00844_ : chn_lut_out_rsci_d_81_70;
  assign _00307_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _03257_ : chn_lut_out_rsci_d_104_82;
  assign _00308_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _00845_ : chn_lut_out_rsci_d_116_105;
  assign _00310_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _03258_ : chn_lut_out_rsci_d_139_117;
  assign _00311_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) lut_in_data_sva_158 : chn_lut_out_rsci_d_267_140;
  assign _00312_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _01775_ : chn_lut_out_rsci_d_268;
  assign _00313_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _01776_ : chn_lut_out_rsci_d_269;
  assign _00314_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _01777_ : chn_lut_out_rsci_d_270;
  assign _00315_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _01778_ : chn_lut_out_rsci_d_271;
  assign _00324_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _03303_ : chn_lut_out_rsci_d_285_280;
  assign _00328_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _03304_ : chn_lut_out_rsci_d_294_289;
  assign _00332_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _03305_ : chn_lut_out_rsci_d_303_298;
  assign _00336_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _03306_ : chn_lut_out_rsci_d_312_307;
  assign _00340_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _02538_ : chn_lut_out_rsci_d_316;
  assign _00341_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _02539_ : chn_lut_out_rsci_d_317;
  assign _00342_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _02540_ : chn_lut_out_rsci_d_318;
  assign _00343_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _02541_ : chn_lut_out_rsci_d_319;
  assign _00344_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _02542_ : chn_lut_out_rsci_d_320;
  assign _00345_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _02543_ : chn_lut_out_rsci_d_321;
  assign _00346_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _02544_ : chn_lut_out_rsci_d_322;
  assign _00347_ = chn_lut_out_and_cse ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7926" *) _02545_ : chn_lut_out_rsci_d_323;
  assign _00306_ = _01774_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7894" *) chn_lut_in_rsci_ld_core_psct_mx0c0 : chn_lut_in_rsci_ld_core_psct;
  assign _00305_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7885" *) _02537_ : chn_lut_in_rsci_iswt0;
  assign _00352_ = core_wen ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7885" *) and_dcpl_72 : chn_lut_out_rsci_iswt0;
  assign nl_lut_lookup_else_1_lo_index_u_1_sva_3 = lut_in_data_sva_154[31:0] - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12655" *) cfg_lut_lo_start_1_sva_41;
  assign nl_lut_lookup_else_1_lo_index_u_2_sva_3 = lut_in_data_sva_154[63:32] - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12665" *) cfg_lut_lo_start_1_sva_41;
  assign nl_lut_lookup_else_1_lo_index_u_3_sva_3[31:0] = lut_in_data_sva_154[95:64] - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12676" *) cfg_lut_lo_start_1_sva_41;
  assign nl_lut_lookup_else_1_lo_index_u_sva_3[31:0] = lut_in_data_sva_154[127:96] - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:12686" *) cfg_lut_lo_start_1_sva_41;
  assign lut_lookup_1_if_else_else_acc_nl = { reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5], _00062_[4:0] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6194" *) { cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5 };
  assign lut_lookup_2_if_else_else_acc_nl = { reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5], _00063_[4:0] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6234" *) { cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5 };
  assign lut_lookup_3_if_else_else_acc_nl = { reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5], _00064_[4:0] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6274" *) { cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5 };
  assign lut_lookup_4_if_else_else_acc_nl = { reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5], _00065_[4:0] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6314" *) { cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5 };
  assign lut_lookup_1_else_1_acc_nl = { cfg_lut_lo_start_rsci_d[31], cfg_lut_lo_start_rsci_d } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6442" *) { chn_lut_in_rsci_d_mxwt[31], chn_lut_in_rsci_d_mxwt[31:0] };
  assign lut_lookup_2_else_1_acc_nl = { cfg_lut_lo_start_rsci_d[31], cfg_lut_lo_start_rsci_d } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6447" *) { chn_lut_in_rsci_d_mxwt[63], chn_lut_in_rsci_d_mxwt[63:32] };
  assign lut_lookup_3_else_1_acc_nl = { cfg_lut_lo_start_rsci_d[31], cfg_lut_lo_start_rsci_d } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6452" *) { chn_lut_in_rsci_d_mxwt[95], chn_lut_in_rsci_d_mxwt[95:64] };
  assign lut_lookup_4_else_1_acc_nl = { cfg_lut_lo_start_rsci_d[31], cfg_lut_lo_start_rsci_d } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6457" *) { chn_lut_in_rsci_d_mxwt[127], chn_lut_in_rsci_d_mxwt[127:96] };
  assign lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0 = lut_in_data_sva_154[31:0] - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6463" *) cfg_lut_le_start_1_sva_41;
  assign lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0 = lut_in_data_sva_154[63:32] - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6466" *) cfg_lut_le_start_1_sva_41;
  assign lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0 = lut_in_data_sva_154[95:64] - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6469" *) cfg_lut_le_start_1_sva_41;
  assign lut_lookup_if_else_else_le_data_sub_sva_mx0w0 = lut_in_data_sva_154[127:96] - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6472" *) cfg_lut_le_start_1_sva_41;
  assign lut_lookup_1_if_if_else_acc_nl = { reg_lut_lookup_1_else_else_else_else_acc_reg, reg_lut_lookup_1_else_else_else_else_acc_reg, reg_lut_lookup_1_else_else_else_else_acc_1_reg, reg_lut_lookup_1_else_else_else_else_acc_2_reg, reg_lut_lookup_1_else_else_else_else_acc_3_reg } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6794" *) { cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7 };
  assign lut_lookup_2_if_if_else_acc_nl = { reg_lut_lookup_2_else_else_else_else_acc_reg, reg_lut_lookup_2_else_else_else_else_acc_reg, reg_lut_lookup_2_else_else_else_else_acc_1_reg, reg_lut_lookup_2_else_else_else_else_acc_2_reg, reg_lut_lookup_2_else_else_else_else_acc_3_reg } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6806" *) { cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7 };
  assign lut_lookup_3_if_if_else_acc_nl = { reg_lut_lookup_3_else_else_else_else_acc_reg, reg_lut_lookup_3_else_else_else_else_acc_reg, reg_lut_lookup_3_else_else_else_else_acc_1_reg, reg_lut_lookup_3_else_else_else_else_acc_2_reg, reg_lut_lookup_3_else_else_else_else_acc_3_reg } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6818" *) { cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7 };
  assign lut_lookup_4_if_if_else_acc_nl = { reg_lut_lookup_4_else_else_else_else_acc_reg, reg_lut_lookup_4_else_else_else_else_acc_reg, reg_lut_lookup_4_else_else_else_else_acc_1_reg, reg_lut_lookup_4_else_else_else_else_acc_2_reg, reg_lut_lookup_4_else_else_else_else_acc_3_reg } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:6830" *) { cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7 };
  assign lut_lookup_if_else_else_else_le_index_s_1_sva = { reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5], _00062_[4:0] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7222" *) { cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5 };
  assign lut_lookup_if_else_else_else_le_index_s_2_sva = { reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5], _00063_[4:0] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7239" *) { cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5 };
  assign lut_lookup_if_else_else_else_le_index_s_3_sva = { reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5], _00064_[4:0] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7256" *) { cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5 };
  assign lut_lookup_if_else_else_else_le_index_s_sva = { reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5], _00065_[4:0] } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7273" *) { cfg_lut_le_index_offset_1_sva_5[7], cfg_lut_le_index_offset_1_sva_5 };
  assign lut_lookup_if_if_else_else_le_index_s_1_sva = { reg_lut_lookup_1_else_else_else_else_acc_reg, reg_lut_lookup_1_else_else_else_else_acc_1_reg, reg_lut_lookup_1_else_else_else_else_acc_2_reg, reg_lut_lookup_1_else_else_else_else_acc_3_reg } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7291" *) { cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7 };
  assign lut_lookup_if_if_else_else_le_index_s_2_sva = { reg_lut_lookup_2_else_else_else_else_acc_reg, reg_lut_lookup_2_else_else_else_else_acc_1_reg, reg_lut_lookup_2_else_else_else_else_acc_2_reg, reg_lut_lookup_2_else_else_else_else_acc_3_reg } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7299" *) { cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7 };
  assign lut_lookup_if_if_else_else_le_index_s_3_sva = { reg_lut_lookup_3_else_else_else_else_acc_reg, reg_lut_lookup_3_else_else_else_else_acc_1_reg, reg_lut_lookup_3_else_else_else_else_acc_2_reg, reg_lut_lookup_3_else_else_else_else_acc_3_reg } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7307" *) { cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7 };
  assign lut_lookup_if_if_else_else_le_index_s_sva = { reg_lut_lookup_4_else_else_else_else_acc_reg, reg_lut_lookup_4_else_else_else_else_acc_1_reg, reg_lut_lookup_4_else_else_else_else_acc_2_reg, reg_lut_lookup_4_else_else_else_else_acc_3_reg } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7315" *) { cfg_lut_le_index_offset_1_sva_7[7], cfg_lut_le_index_offset_1_sva_7 };
  assign lut_lookup_1_else_else_acc_1_nl = { cfg_lut_le_start_rsci_d[31], cfg_lut_le_start_rsci_d } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7318" *) { chn_lut_in_rsci_d_mxwt[31], chn_lut_in_rsci_d_mxwt[31:0] };
  assign lut_lookup_3_else_else_acc_1_nl = { cfg_lut_le_start_rsci_d[31], cfg_lut_le_start_rsci_d } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7322" *) { chn_lut_in_rsci_d_mxwt[95], chn_lut_in_rsci_d_mxwt[95:64] };
  assign lut_lookup_2_else_else_acc_1_nl = { cfg_lut_le_start_rsci_d[31], cfg_lut_le_start_rsci_d } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7328" *) { chn_lut_in_rsci_d_mxwt[63], chn_lut_in_rsci_d_mxwt[63:32] };
  assign lut_lookup_4_else_else_acc_1_nl = { cfg_lut_le_start_rsci_d[31], cfg_lut_le_start_rsci_d } - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:7333" *) { chn_lut_in_rsci_d_mxwt[127], chn_lut_in_rsci_d_mxwt[127:96] };
  assign _03905_ = and_896_cse ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5989" *) cfg_lut_le_function_1_sva_st_41;
  assign _03906_ = chn_lut_in_rsci_d_mxwt[31] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8141" *) cfg_lut_le_start_rsci_d[31];
  assign _03907_ = chn_lut_in_rsci_d_mxwt[31] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8155" *) cfg_lut_lo_start_rsci_d[31];
  assign _03908_ = chn_lut_in_rsci_d_mxwt[63] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8192" *) cfg_lut_le_start_rsci_d[31];
  assign _03909_ = chn_lut_in_rsci_d_mxwt[63] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8194" *) cfg_lut_lo_start_rsci_d[31];
  assign _03910_ = chn_lut_in_rsci_d_mxwt[95] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8196" *) cfg_lut_le_start_rsci_d[31];
  assign _03911_ = chn_lut_in_rsci_d_mxwt[95] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8199" *) cfg_lut_lo_start_rsci_d[31];
  assign _03912_ = chn_lut_in_rsci_d_mxwt[127] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8202" *) cfg_lut_le_start_rsci_d[31];
  assign _03913_ = chn_lut_in_rsci_d_mxwt[127] ^ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:8204" *) cfg_lut_lo_start_rsci_d[31];
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5404" *)
  NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_in_rsci_inst (
    .chn_lut_in_rsc_lz(chn_lut_in_rsc_lz),
    .chn_lut_in_rsc_vz(chn_lut_in_rsc_vz),
    .chn_lut_in_rsc_z(chn_lut_in_rsc_z),
    .chn_lut_in_rsci_bawt(chn_lut_in_rsci_bawt),
    .chn_lut_in_rsci_d_mxwt(chn_lut_in_rsci_d_mxwt),
    .chn_lut_in_rsci_iswt0(chn_lut_in_rsci_iswt0),
    .chn_lut_in_rsci_ld_core_psct(chn_lut_in_rsci_ld_core_psct),
    .chn_lut_in_rsci_oswt(chn_lut_in_rsci_oswt),
    .chn_lut_in_rsci_wen_comp(chn_lut_in_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5420" *)
  NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_inst (
    .chn_lut_out_rsc_lz(chn_lut_out_rsc_lz),
    .chn_lut_out_rsc_vz(chn_lut_out_rsc_vz),
    .chn_lut_out_rsc_z(chn_lut_out_rsc_z),
    .chn_lut_out_rsci_bawt(chn_lut_out_rsci_bawt),
    .chn_lut_out_rsci_d({ chn_lut_out_rsci_d_323, chn_lut_out_rsci_d_322, chn_lut_out_rsci_d_321, chn_lut_out_rsci_d_320, chn_lut_out_rsci_d_319, chn_lut_out_rsci_d_318, chn_lut_out_rsci_d_317, chn_lut_out_rsci_d_316, chn_lut_out_rsci_d_315, chn_lut_out_rsci_d_314, chn_lut_out_rsci_d_313, chn_lut_out_rsci_d_312_307, chn_lut_out_rsci_d_306, chn_lut_out_rsci_d_305, chn_lut_out_rsci_d_304, chn_lut_out_rsci_d_303_298, chn_lut_out_rsci_d_297, chn_lut_out_rsci_d_296, chn_lut_out_rsci_d_295, chn_lut_out_rsci_d_294_289, chn_lut_out_rsci_d_288, chn_lut_out_rsci_d_287, chn_lut_out_rsci_d_286, chn_lut_out_rsci_d_285_280, chn_lut_out_rsci_d_279, chn_lut_out_rsci_d_278, chn_lut_out_rsci_d_277, chn_lut_out_rsci_d_276, chn_lut_out_rsci_d_275, chn_lut_out_rsci_d_274, chn_lut_out_rsci_d_273, chn_lut_out_rsci_d_272, chn_lut_out_rsci_d_271, chn_lut_out_rsci_d_270, chn_lut_out_rsci_d_269, chn_lut_out_rsci_d_268, chn_lut_out_rsci_d_267_140, chn_lut_out_rsci_d_139_117, chn_lut_out_rsci_d_116_105, chn_lut_out_rsci_d_104_82, chn_lut_out_rsci_d_81_70, chn_lut_out_rsci_d_69_47, chn_lut_out_rsci_d_46_35, chn_lut_out_rsci_d_34_12, chn_lut_out_rsci_d_11_0 }),
    .chn_lut_out_rsci_iswt0(chn_lut_out_rsci_iswt0),
    .chn_lut_out_rsci_ld_core_psct(reg_chn_lut_out_rsci_ld_core_psct_cse),
    .chn_lut_out_rsci_oswt(chn_lut_out_rsci_oswt),
    .chn_lut_out_rsci_wen_comp(chn_lut_out_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5445" *)
  NV_NVDLA_SDP_CORE_Y_idx_core_core_fsm NV_NVDLA_SDP_CORE_Y_idx_core_core_fsm_inst (
    .core_wen(core_wen),
    .fsm_output(fsm_output),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5436" *)
  NV_NVDLA_SDP_CORE_Y_idx_core_staller NV_NVDLA_SDP_CORE_Y_idx_core_staller_inst (
    .chn_lut_in_rsci_wen_comp(chn_lut_in_rsci_wen_comp),
    .chn_lut_out_rsci_wen_comp(chn_lut_out_rsci_wen_comp),
    .core_wen(core_wen),
    .core_wten(core_wten),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4698" *)
  \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=10\width=1  cfg_lut_hybrid_priority_rsci (
    .d(cfg_lut_hybrid_priority_rsci_d),
    .z(cfg_lut_hybrid_priority_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4683" *)
  \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=7\width=1  cfg_lut_le_function_rsci (
    .d(cfg_lut_le_function_rsci_d),
    .z(cfg_lut_le_function_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4668" *)
  \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=4\width=8  cfg_lut_le_index_offset_rsci (
    .d(cfg_lut_le_index_offset_rsci_d),
    .z(cfg_lut_le_index_offset_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4673" *)
  \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=5\width=8  cfg_lut_le_index_select_rsci (
    .d(cfg_lut_le_index_select_rsci_d),
    .z(cfg_lut_le_index_select_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4658" *)
  \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=2\width=32  cfg_lut_le_start_rsci (
    .d(cfg_lut_le_start_rsci_d),
    .z(cfg_lut_le_start_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4678" *)
  \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=6\width=8  cfg_lut_lo_index_select_rsci (
    .d(cfg_lut_lo_index_select_rsci_d),
    .z(cfg_lut_lo_index_select_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4663" *)
  \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=3\width=32  cfg_lut_lo_start_rsci (
    .d(cfg_lut_lo_start_rsci_d),
    .z(cfg_lut_lo_start_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4693" *)
  \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=9\width=1  cfg_lut_oflow_priority_rsci (
    .d(cfg_lut_oflow_priority_rsci_d),
    .z(cfg_lut_oflow_priority_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4688" *)
  \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=8\width=1  cfg_lut_uflow_priority_rsci (
    .d(cfg_lut_uflow_priority_rsci_d),
    .z(cfg_lut_uflow_priority_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4703" *)
  \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=11\width=2  cfg_precision_rsci (
    .d(cfg_precision_rsci_d),
    .z(cfg_precision_rsc_z)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5084" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, lut_in_data_sva_154[22:0] }),
    .s({ lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_1_a_int_mant_p1_1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5076" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] }),
    .s({ lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5100" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_1_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2, lut_in_data_sva_154[22:0] }),
    .s({ lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl, nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_2_a_int_mant_p1_1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5092" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2, cfg_lut_lo_start_1_sva_41[22:0] }),
    .s({ _02029_[7:4], lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl, nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_2_addend_larger_asn_19_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5068" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, lut_in_data_sva_154[22:0] }),
    .s({ lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_a_int_mant_p1_1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5060" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] }),
    .s({ lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_addend_larger_asn_19_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4742" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=35  lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg (
    .a({ 1'b1, FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5 }),
    .s(nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s),
    .z(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4751" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=10\width_z=256  lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg (
    .a({ 1'b1, FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5 }),
    .s(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp),
    .z(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4724" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=35  lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg (
    .a({ 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm }),
    .s(nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s[8:0]),
    .z(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4733" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=10\width_z=256  lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg (
    .a({ 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm }),
    .s(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp),
    .z(lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5269" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_rg (
    .a(FpAdd_8U_23U_2_int_mant_p1_1_sva_3[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13),
    .z(lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5252" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  lut_lookup_1_FpNormalize_8U_49U_else_lshift_rg (
    .a(FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12),
    .z(lut_lookup_1_FpNormalize_8U_49U_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4996" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=32\width_z=31  lut_lookup_1_IntLog2_32U_lshift_rg (
    .a(1'b1),
    .s({ reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], nl_lut_lookup_1_IntLog2_32U_lshift_rg_s[4:0] }),
    .z(lut_lookup_1_IntLog2_32U_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5277" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=159\signd_a=0\width_s=8\width_z=287  lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg (
    .a({ lut_lookup_else_1_lo_index_u_1_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_lut_lo_index_select_1_sva_5),
    .z(lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5260" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=159\signd_a=0\width_s=8\width_z=287  lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg (
    .a({ lut_lookup_else_else_else_le_index_u_1_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_lut_le_index_select_1_sva_5),
    .z(lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5396" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=1\signd_a=0\width_s=8\width_z=32  lut_lookup_1_else_1_else_else_lo_data_f_lshift_1_rg (
    .a(1'b1),
    .s(cfg_lut_lo_index_select_1_sva_6),
    .z(lut_lookup_1_else_1_else_else_lo_data_f_lshift_1_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4892" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=32\signd_a=0\width_s=9\width_z=35  lut_lookup_1_else_1_else_else_rshift_rg (
    .a(lut_lookup_1_else_1_else_else_lo_data_f_and_itm_2),
    .s({ reg_lut_lookup_1_else_1_else_else_acc_itm, reg_lut_lookup_1_else_1_else_else_acc_1_itm }),
    .z(lut_lookup_1_else_1_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5388" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=1\signd_a=0\width_s=8\width_z=32  lut_lookup_1_else_else_else_else_le_data_f_lshift_1_rg (
    .a(1'b1),
    .s(cfg_lut_le_index_select_1_sva_6),
    .z(lut_lookup_1_else_else_else_else_le_data_f_lshift_1_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4884" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=35\signd_a=0\width_s=9\width_z=35  lut_lookup_1_else_else_else_else_rshift_rg (
    .a({ lut_lookup_1_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_1_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_1_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_1_else_else_else_else_le_data_f_and_itm_2 }),
    .s({ reg_lut_lookup_1_else_else_else_else_acc_reg, reg_lut_lookup_1_else_else_else_else_acc_1_reg, reg_lut_lookup_1_else_else_else_else_acc_2_reg, reg_lut_lookup_1_else_else_else_else_acc_3_reg }),
    .z(lut_lookup_1_else_else_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4876" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=31\signd_a=0\width_s=8\width_z=35  lut_lookup_1_if_else_else_else_else_else_rshift_rg (
    .a({ reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm, reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm }),
    .s({ 1'b1, reg_lut_lookup_1_else_else_else_else_acc_2_reg, reg_lut_lookup_1_else_else_else_else_acc_3_reg }),
    .z(lut_lookup_1_if_else_else_else_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4868" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=31\signd_a=0\width_s=6\width_z=35  lut_lookup_1_if_else_else_else_else_if_lshift_rg (
    .a({ reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm, reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm }),
    .s({ reg_lut_lookup_1_else_else_else_else_acc_3_reg, lut_lookup_1_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 }),
    .z(lut_lookup_1_if_else_else_else_else_if_lshift_itm)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4708" *)
  SDP_Y_IDX_leading_sign_32_0 lut_lookup_1_leading_sign_32_0_rg (
    .mantissa(lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0),
    .rtn(libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_4)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5032" *)
  SDP_Y_IDX_leading_sign_49_0 lut_lookup_1_leading_sign_49_0_2_rg (
    .mantissa(FpAdd_8U_23U_2_int_mant_p1_1_sva_3[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5028" *)
  SDP_Y_IDX_leading_sign_49_0 lut_lookup_1_leading_sign_49_0_rg (
    .mantissa(FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5132" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, lut_in_data_sva_154[54:32] }),
    .s({ lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_1_a_int_mant_p1_2_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5124" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] }),
    .s({ lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5148" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_2_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2, lut_in_data_sva_154[54:32] }),
    .s({ lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl, nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_2_a_int_mant_p1_2_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5140" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2, cfg_lut_lo_start_1_sva_41[22:0] }),
    .s({ lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl, nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_2_addend_larger_asn_13_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5116" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, lut_in_data_sva_154[54:32] }),
    .s({ lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_a_int_mant_p1_2_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5108" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] }),
    .s({ lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_addend_larger_asn_13_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4778" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=35  lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg (
    .a({ 1'b1, FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5 }),
    .s(nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s),
    .z(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4787" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=10\width_z=256  lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg (
    .a({ 1'b1, FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5 }),
    .s(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp),
    .z(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4760" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=35  lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg (
    .a({ 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg }),
    .s(nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s[8:0]),
    .z(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4769" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=10\width_z=256  lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg (
    .a({ 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg }),
    .s(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp),
    .z(lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5303" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_rg (
    .a(FpAdd_8U_23U_2_int_mant_p1_2_sva_3[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15),
    .z(lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5286" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  lut_lookup_2_FpNormalize_8U_49U_else_lshift_rg (
    .a(FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14),
    .z(lut_lookup_2_FpNormalize_8U_49U_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5004" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=32\width_z=31  lut_lookup_2_IntLog2_32U_lshift_rg (
    .a(1'b1),
    .s({ reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], nl_lut_lookup_2_IntLog2_32U_lshift_rg_s[4:0] }),
    .z(lut_lookup_2_IntLog2_32U_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5311" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=159\signd_a=0\width_s=8\width_z=287  lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg (
    .a({ lut_lookup_else_1_lo_index_u_2_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_lut_lo_index_select_1_sva_5),
    .z(lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5294" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=159\signd_a=0\width_s=8\width_z=287  lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg (
    .a({ lut_lookup_else_else_else_le_index_u_2_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_lut_le_index_select_1_sva_5),
    .z(lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4924" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=32\signd_a=0\width_s=9\width_z=35  lut_lookup_2_else_1_else_else_rshift_rg (
    .a(lut_lookup_2_else_1_else_else_lo_data_f_and_itm_2),
    .s({ reg_lut_lookup_2_else_1_else_else_acc_itm, reg_lut_lookup_2_else_1_else_else_acc_1_itm }),
    .z(lut_lookup_2_else_1_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4916" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=35\signd_a=0\width_s=9\width_z=35  lut_lookup_2_else_else_else_else_rshift_rg (
    .a({ lut_lookup_2_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_2_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_2_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_2_else_else_else_else_le_data_f_and_itm_2 }),
    .s({ reg_lut_lookup_2_else_else_else_else_acc_reg, reg_lut_lookup_2_else_else_else_else_acc_1_reg, reg_lut_lookup_2_else_else_else_else_acc_2_reg, reg_lut_lookup_2_else_else_else_else_acc_3_reg }),
    .z(lut_lookup_2_else_else_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4908" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=31\signd_a=0\width_s=8\width_z=35  lut_lookup_2_if_else_else_else_else_else_rshift_rg (
    .a({ reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg }),
    .s({ 1'b1, reg_lut_lookup_2_else_else_else_else_acc_2_reg, reg_lut_lookup_2_else_else_else_else_acc_3_reg }),
    .z(lut_lookup_2_if_else_else_else_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4900" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=31\signd_a=0\width_s=6\width_z=35  lut_lookup_2_if_else_else_else_else_if_lshift_rg (
    .a({ reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg }),
    .s({ reg_lut_lookup_2_else_else_else_else_acc_3_reg, lut_lookup_2_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 }),
    .z(lut_lookup_2_if_else_else_else_else_if_lshift_itm)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4712" *)
  SDP_Y_IDX_leading_sign_32_0 lut_lookup_2_leading_sign_32_0_rg (
    .mantissa(lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0),
    .rtn(libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_5)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5040" *)
  SDP_Y_IDX_leading_sign_49_0 lut_lookup_2_leading_sign_49_0_2_rg (
    .mantissa(FpAdd_8U_23U_2_int_mant_p1_2_sva_3[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5036" *)
  SDP_Y_IDX_leading_sign_49_0 lut_lookup_2_leading_sign_49_0_rg (
    .mantissa(FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5180" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, lut_in_data_sva_154[86:64] }),
    .s({ lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_1_a_int_mant_p1_3_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5172" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] }),
    .s({ lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5196" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_3_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2, lut_in_data_sva_154[86:64] }),
    .s({ lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl, nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_2_a_int_mant_p1_3_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5188" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2, cfg_lut_lo_start_1_sva_41[22:0] }),
    .s({ lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl, nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_2_addend_larger_asn_7_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5164" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, lut_in_data_sva_154[86:64] }),
    .s({ lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_a_int_mant_p1_3_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5156" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] }),
    .s({ lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_addend_larger_asn_7_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4814" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=35  lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg (
    .a({ 1'b1, FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5 }),
    .s(nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s),
    .z(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4823" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=10\width_z=256  lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg (
    .a({ 1'b1, FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5 }),
    .s(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp),
    .z(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4796" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=35  lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg (
    .a({ 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg }),
    .s(nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s[8:0]),
    .z(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4805" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=10\width_z=256  lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg (
    .a({ 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg }),
    .s(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp),
    .z(lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5337" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_rg (
    .a(FpAdd_8U_23U_2_int_mant_p1_3_sva_3[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_17),
    .z(lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5320" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  lut_lookup_3_FpNormalize_8U_49U_else_lshift_rg (
    .a(FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_16),
    .z(lut_lookup_3_FpNormalize_8U_49U_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5012" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=32\width_z=31  lut_lookup_3_IntLog2_32U_lshift_rg (
    .a(1'b1),
    .s({ reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], nl_lut_lookup_3_IntLog2_32U_lshift_rg_s[4:0] }),
    .z(lut_lookup_3_IntLog2_32U_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5345" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=159\signd_a=0\width_s=8\width_z=287  lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg (
    .a({ lut_lookup_else_1_lo_index_u_3_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_lut_lo_index_select_1_sva_5),
    .z(lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5328" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=159\signd_a=0\width_s=8\width_z=287  lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg (
    .a({ lut_lookup_else_else_else_le_index_u_3_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_lut_le_index_select_1_sva_5),
    .z(lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4956" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=32\signd_a=0\width_s=9\width_z=35  lut_lookup_3_else_1_else_else_rshift_rg (
    .a(lut_lookup_3_else_1_else_else_lo_data_f_and_itm_2),
    .s({ reg_lut_lookup_3_else_1_else_else_acc_itm, reg_lut_lookup_3_else_1_else_else_acc_1_itm }),
    .z(lut_lookup_3_else_1_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4948" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=35\signd_a=0\width_s=9\width_z=35  lut_lookup_3_else_else_else_else_rshift_rg (
    .a({ lut_lookup_3_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_3_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_3_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_3_else_else_else_else_le_data_f_and_itm_2 }),
    .s({ reg_lut_lookup_3_else_else_else_else_acc_reg, reg_lut_lookup_3_else_else_else_else_acc_1_reg, reg_lut_lookup_3_else_else_else_else_acc_2_reg, reg_lut_lookup_3_else_else_else_else_acc_3_reg }),
    .z(lut_lookup_3_else_else_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4940" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=31\signd_a=0\width_s=8\width_z=35  lut_lookup_3_if_else_else_else_else_else_rshift_rg (
    .a({ reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg }),
    .s({ 1'b1, reg_lut_lookup_3_else_else_else_else_acc_2_reg, reg_lut_lookup_3_else_else_else_else_acc_3_reg }),
    .z(lut_lookup_3_if_else_else_else_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4932" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=31\signd_a=0\width_s=6\width_z=35  lut_lookup_3_if_else_else_else_else_if_lshift_rg (
    .a({ reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg }),
    .s({ reg_lut_lookup_3_else_else_else_else_acc_3_reg, lut_lookup_3_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 }),
    .z(lut_lookup_3_if_else_else_else_else_if_lshift_itm)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4716" *)
  SDP_Y_IDX_leading_sign_32_0 lut_lookup_3_leading_sign_32_0_rg (
    .mantissa(lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0),
    .rtn(libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_6)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5048" *)
  SDP_Y_IDX_leading_sign_49_0 lut_lookup_3_leading_sign_49_0_2_rg (
    .mantissa(FpAdd_8U_23U_2_int_mant_p1_3_sva_3[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_17)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5044" *)
  SDP_Y_IDX_leading_sign_49_0 lut_lookup_3_leading_sign_49_0_rg (
    .mantissa(FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_16)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5228" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, lut_in_data_sva_154[118:96] }),
    .s({ lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_1_a_int_mant_p1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5220" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] }),
    .s({ lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5244" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2, lut_in_data_sva_154[118:96] }),
    .s({ lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl, nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_2_a_int_mant_p1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5236" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2, cfg_lut_lo_start_1_sva_41[22:0] }),
    .s({ lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl, nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_2_addend_larger_asn_1_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5212" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
    .a({ lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, lut_in_data_sva_154[118:96] }),
    .s({ lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_a_int_mant_p1_sva)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5204" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=49  lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
    .a({ lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] }),
    .s({ lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] }),
    .z(FpAdd_8U_23U_addend_larger_asn_1_mx0w1)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4850" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=35  lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg (
    .a({ 1'b1, FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5 }),
    .s(nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_s),
    .z(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4859" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=10\width_z=256  lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg (
    .a({ 1'b1, FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5 }),
    .s(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp),
    .z(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4832" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=9\width_z=35  lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg (
    .a({ 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 }),
    .s({ _02030_[8], nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s }),
    .z(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4841" *)
  \$paramod\SDP_Y_IDX_mgc_shift_bl_v4\width_a=24\signd_a=0\width_s=10\width_z=256  lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg (
    .a({ 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 }),
    .s(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp),
    .z(lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5371" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_rg (
    .a(FpAdd_8U_23U_2_int_mant_p1_sva_3[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_19),
    .z(lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5354" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=49\signd_a=0\width_s=6\width_z=49  lut_lookup_4_FpNormalize_8U_49U_else_lshift_rg (
    .a(FpAdd_8U_23U_1_int_mant_p1_sva_3[48:0]),
    .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_18),
    .z(lut_lookup_4_FpNormalize_8U_49U_else_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5020" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=1\signd_a=0\width_s=32\width_z=31  lut_lookup_4_IntLog2_32U_lshift_rg (
    .a(1'b1),
    .s({ reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], nl_lut_lookup_4_IntLog2_32U_lshift_rg_s[4:0] }),
    .z(lut_lookup_4_IntLog2_32U_lshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5379" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=159\signd_a=0\width_s=8\width_z=287  lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg (
    .a({ lut_lookup_else_1_lo_index_u_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_lut_lo_index_select_1_sva_5),
    .z(lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5362" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=159\signd_a=0\width_s=8\width_z=287  lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg (
    .a({ lut_lookup_else_else_else_le_index_u_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 }),
    .s(cfg_lut_le_index_select_1_sva_5),
    .z(lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4988" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=32\signd_a=0\width_s=9\width_z=35  lut_lookup_4_else_1_else_else_rshift_rg (
    .a(lut_lookup_4_else_1_else_else_lo_data_f_and_itm_2),
    .s({ reg_lut_lookup_4_else_1_else_else_acc_itm, reg_lut_lookup_4_else_1_else_else_acc_1_itm }),
    .z(lut_lookup_4_else_1_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4980" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=35\signd_a=0\width_s=9\width_z=35  lut_lookup_4_else_else_else_else_rshift_rg (
    .a({ lut_lookup_4_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_4_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_4_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_4_else_else_else_else_le_data_f_and_itm_2 }),
    .s({ reg_lut_lookup_4_else_else_else_else_acc_reg, reg_lut_lookup_4_else_else_else_else_acc_1_reg, reg_lut_lookup_4_else_else_else_else_acc_2_reg, reg_lut_lookup_4_else_else_else_else_acc_3_reg }),
    .z(lut_lookup_4_else_else_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4972" *)
  \$paramod\SDP_Y_IDX_mgc_shift_br_v4\width_a=31\signd_a=0\width_s=8\width_z=35  lut_lookup_4_if_else_else_else_else_else_rshift_rg (
    .a({ reg_IntLog2_32U_ac_int_cctor_1_30_0_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 }),
    .s({ 1'b1, reg_lut_lookup_4_else_else_else_else_acc_2_reg, reg_lut_lookup_4_else_else_else_else_acc_3_reg }),
    .z(lut_lookup_4_if_else_else_else_else_else_rshift_itm)
  );
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4964" *)
  \$paramod\SDP_Y_IDX_mgc_shift_l_v4\width_a=31\signd_a=0\width_s=6\width_z=35  lut_lookup_4_if_else_else_else_else_if_lshift_rg (
    .a({ reg_IntLog2_32U_ac_int_cctor_1_30_0_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 }),
    .s({ reg_lut_lookup_4_else_else_else_else_acc_3_reg, lut_lookup_4_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 }),
    .z(lut_lookup_4_if_else_else_else_else_if_lshift_itm)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:4720" *)
  SDP_Y_IDX_leading_sign_32_0 lut_lookup_4_leading_sign_32_0_rg (
    .mantissa(lut_lookup_if_else_else_le_data_sub_sva_mx0w0),
    .rtn(libraries_leading_sign_32_0_bddfe7269a66a92265caaec08a257f83661f_7)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5056" *)
  SDP_Y_IDX_leading_sign_49_0 lut_lookup_4_leading_sign_49_0_2_rg (
    .mantissa(FpAdd_8U_23U_2_int_mant_p1_sva_3[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_19)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:5052" *)
  SDP_Y_IDX_leading_sign_49_0 lut_lookup_4_leading_sign_49_0_rg (
    .mantissa(FpAdd_8U_23U_1_int_mant_p1_sva_3[48:0]),
    .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_18)
  );
  assign _00062_[8:5] = { reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_2_lpi_1_dfm_4_1_itm[5] };
  assign _00063_[8:5] = { reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_3_lpi_1_dfm_4_1_itm[5] };
  assign _00064_[8:5] = { reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_4_lpi_1_dfm_4_1_itm[5] };
  assign _00065_[8:5] = { reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5], reg_FpAdd_8U_23U_1_qr_lpi_1_dfm_4_1_itm[5] };
  assign _00066_[6] = _00066_[7];
  assign _00067_[6] = _00067_[7];
  assign _00070_[33:0] = { _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34], _00070_[34] };
  assign _00071_[33:0] = { _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34], _00071_[34] };
  assign _00072_[33:0] = { _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34], _00072_[34] };
  assign _00073_[33:0] = { _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34], _00073_[34] };
  assign _00074_[33:0] = { _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34], _00074_[34] };
  assign _00075_[33:0] = { _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34], _00075_[34] };
  assign _00076_[33:0] = { _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34], _00076_[34] };
  assign _00077_[33:0] = { _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34], _00077_[34] };
  assign _00078_[33:0] = { _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34], _00078_[34] };
  assign _00079_[33:0] = { _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34], _00079_[34] };
  assign _00080_[33:0] = { _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34], _00080_[34] };
  assign _00081_[33:0] = { _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34], _00081_[34] };
  assign _00082_[33:0] = { _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34], _00082_[34] };
  assign _00083_[33:0] = { _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34], _00083_[34] };
  assign _00084_[33:0] = { _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34], _00084_[34] };
  assign _00085_[33:0] = { _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34], _00085_[34] };
  assign _00086_[33:0] = { _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34], _00086_[34] };
  assign _00087_[33:0] = { _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34], _00087_[34] };
  assign _00088_[33:0] = { _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34], _00088_[34] };
  assign _00089_[33:0] = { _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34], _00089_[34] };
  assign _02027_[5:0] = _01007_;
  assign _02029_[3:0] = lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  assign _02030_[7:0] = nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_s;
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_cse = FpMantRNE_49U_24U_2_else_carry_FpMantRNE_49U_24U_2_else_carry_or_3_cse;
  assign FpAdd_8U_23U_1_is_a_greater_acc_10_itm_8_1 = FpAdd_8U_23U_1_is_a_greater_acc_10_nl[8];
  assign FpAdd_8U_23U_1_is_a_greater_acc_4_itm_8_1 = FpAdd_8U_23U_1_is_a_greater_acc_4_nl[8];
  assign FpAdd_8U_23U_1_is_a_greater_acc_6_itm_8_1 = FpAdd_8U_23U_1_is_a_greater_acc_6_nl[8];
  assign FpAdd_8U_23U_1_is_a_greater_acc_8_itm_8_1 = FpAdd_8U_23U_1_is_a_greater_acc_8_nl[8];
  assign FpAdd_8U_23U_1_is_inf_and_1_cse = FpAdd_8U_23U_2_is_inf_and_cse;
  assign FpAdd_8U_23U_2_is_a_greater_acc_1_itm_8_1 = FpAdd_8U_23U_2_is_a_greater_acc_1_nl[8];
  assign FpAdd_8U_23U_2_is_a_greater_acc_2_itm_8_1 = FpAdd_8U_23U_2_is_a_greater_acc_2_nl[8];
  assign FpAdd_8U_23U_2_is_a_greater_acc_3_itm_8_1 = FpAdd_8U_23U_2_is_a_greater_acc_3_nl[8];
  assign FpAdd_8U_23U_2_is_a_greater_acc_itm_8_1 = FpAdd_8U_23U_2_is_a_greater_acc_nl[8];
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_itm_23_1 = FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl[23];
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_itm_23_1 = FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl[23];
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_itm_23_1 = FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl[23];
  assign FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_itm_23_1 = FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl[23];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_itm_23_1 = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl[23];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_itm_23_1 = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl[23];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_itm_23_1 = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl[23];
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_itm_23_1 = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl[23];
  assign IsNaN_8U_23U_7_aelse_and_17_cse = IsNaN_8U_23U_1_aelse_and_4_cse;
  assign and_574_rgt = and_564_rgt;
  assign and_636_cse = and_428_rgt;
  assign chn_lut_in_rsci_oswt_unreg = or_tmp_1628;
  assign lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 = lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7];
  assign lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1 = lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7];
  assign lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 = lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7];
  assign lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1 = lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7];
  assign lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1 = lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247];
  assign lut_lookup_1_else_1_acc_itm_32 = lut_lookup_1_else_1_acc_nl[32];
  assign lut_lookup_1_else_else_acc_1_itm_32 = lut_lookup_1_else_else_acc_1_nl[32];
  assign lut_lookup_1_else_else_else_if_acc_itm_3_1 = lut_lookup_1_else_else_else_if_acc_nl[3];
  assign lut_lookup_1_else_if_else_if_acc_itm_3_1 = lut_lookup_1_else_if_else_if_acc_nl[3];
  assign lut_lookup_1_if_else_else_acc_itm_10 = lut_lookup_1_if_else_else_acc_nl[10];
  assign lut_lookup_1_if_else_else_else_else_acc_itm_32_1 = lut_lookup_1_if_else_else_else_else_acc_nl[32];
  assign lut_lookup_1_if_else_else_else_if_acc_itm_3 = lut_lookup_1_if_else_else_else_if_acc_nl[3];
  assign lut_lookup_1_if_if_else_acc_itm_9_1 = lut_lookup_1_if_if_else_acc_nl[9];
  assign lut_lookup_1_if_if_else_else_if_acc_itm_3 = lut_lookup_1_if_if_else_else_if_acc_nl[3];
  assign lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 = lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7];
  assign lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1 = lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7];
  assign lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 = lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7];
  assign lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1 = lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7];
  assign lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1 = lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247];
  assign lut_lookup_2_else_1_acc_itm_32 = lut_lookup_2_else_1_acc_nl[32];
  assign lut_lookup_2_else_else_acc_1_itm_32 = lut_lookup_2_else_else_acc_1_nl[32];
  assign lut_lookup_2_else_else_else_if_acc_itm_3_1 = lut_lookup_2_else_else_else_if_acc_nl[3];
  assign lut_lookup_2_else_if_else_if_acc_itm_3_1 = lut_lookup_2_else_if_else_if_acc_nl[3];
  assign lut_lookup_2_if_else_else_acc_itm_10 = lut_lookup_2_if_else_else_acc_nl[10];
  assign lut_lookup_2_if_else_else_else_else_acc_itm_32_1 = lut_lookup_2_if_else_else_else_else_acc_nl[32];
  assign lut_lookup_2_if_else_else_else_if_acc_itm_3_1 = lut_lookup_2_if_else_else_else_if_acc_nl[3];
  assign lut_lookup_2_if_if_else_acc_itm_9_1 = lut_lookup_2_if_if_else_acc_nl[9];
  assign lut_lookup_2_if_if_else_else_if_acc_itm_3 = lut_lookup_2_if_if_else_else_if_acc_nl[3];
  assign lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 = lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7];
  assign lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1 = lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7];
  assign lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 = lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7];
  assign lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1 = lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7];
  assign lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1 = lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247];
  assign lut_lookup_3_else_1_acc_itm_32 = lut_lookup_3_else_1_acc_nl[32];
  assign lut_lookup_3_else_else_acc_1_itm_32 = lut_lookup_3_else_else_acc_1_nl[32];
  assign lut_lookup_3_else_else_else_if_acc_itm_3_1 = lut_lookup_3_else_else_else_if_acc_nl[3];
  assign lut_lookup_3_else_if_else_if_acc_itm_3_1 = lut_lookup_3_else_if_else_if_acc_nl[3];
  assign lut_lookup_3_if_else_else_acc_itm_10 = lut_lookup_3_if_else_else_acc_nl[10];
  assign lut_lookup_3_if_else_else_else_else_acc_itm_32_1 = lut_lookup_3_if_else_else_else_else_acc_nl[32];
  assign lut_lookup_3_if_else_else_else_if_acc_itm_3_1 = lut_lookup_3_if_else_else_else_if_acc_nl[3];
  assign lut_lookup_3_if_if_else_acc_itm_9_1 = lut_lookup_3_if_if_else_acc_nl[9];
  assign lut_lookup_3_if_if_else_else_if_acc_itm_3 = lut_lookup_3_if_if_else_else_if_acc_nl[3];
  assign lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_itm_7 = lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7];
  assign lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_itm_7_1 = lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7];
  assign lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_itm_7_1 = lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7];
  assign lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_itm_7_1 = lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7];
  assign lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_itm_247_1 = lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247];
  assign lut_lookup_4_else_1_acc_itm_32 = lut_lookup_4_else_1_acc_nl[32];
  assign lut_lookup_4_else_else_acc_1_itm_32 = lut_lookup_4_else_else_acc_1_nl[32];
  assign lut_lookup_4_else_else_else_if_acc_itm_3_1 = lut_lookup_4_else_else_else_if_acc_nl[3];
  assign lut_lookup_4_else_if_else_if_acc_itm_3_1 = lut_lookup_4_else_if_else_if_acc_nl[3];
  assign lut_lookup_4_if_else_else_acc_itm_10 = lut_lookup_4_if_else_else_acc_nl[10];
  assign lut_lookup_4_if_else_else_else_else_acc_itm_32_1 = lut_lookup_4_if_else_else_else_else_acc_nl[32];
  assign lut_lookup_4_if_else_else_else_if_acc_itm_3_1 = lut_lookup_4_if_else_else_else_if_acc_nl[3];
  assign lut_lookup_4_if_if_else_acc_itm_9_1 = lut_lookup_4_if_if_else_acc_nl[9];
  assign lut_lookup_4_if_if_else_else_if_acc_itm_3 = lut_lookup_4_if_if_else_else_if_acc_nl[3];
  assign lut_lookup_else_1_lut_lookup_lo_uflow_or_3_cse = lut_lookup_if_else_else_else_else_if_lut_lookup_if_else_else_else_else_if_or_3_cse;
  assign mux_314_nl = mux_272_nl;
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_10_nl[8:0] = FpAdd_8U_23U_1_is_a_greater_acc_10_nl;
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_4_nl[8:0] = FpAdd_8U_23U_1_is_a_greater_acc_4_nl;
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_6_nl[8:0] = FpAdd_8U_23U_1_is_a_greater_acc_6_nl;
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_8_nl[8:0] = FpAdd_8U_23U_1_is_a_greater_acc_8_nl;
  assign nl_FpAdd_8U_23U_2_is_a_greater_acc_1_nl[8:0] = FpAdd_8U_23U_2_is_a_greater_acc_1_nl;
  assign nl_FpAdd_8U_23U_2_is_a_greater_acc_2_nl[8:0] = FpAdd_8U_23U_2_is_a_greater_acc_2_nl;
  assign nl_FpAdd_8U_23U_2_is_a_greater_acc_3_nl[8:0] = FpAdd_8U_23U_2_is_a_greater_acc_3_nl;
  assign nl_FpAdd_8U_23U_2_is_a_greater_acc_nl[8:0] = FpAdd_8U_23U_2_is_a_greater_acc_nl;
  assign nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl[23:0] = FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_1_nl;
  assign nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl[23:0] = FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_2_nl;
  assign nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl[23:0] = FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_3_nl;
  assign nl_FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl[23:0] = FpAdd_8U_23U_2_is_a_greater_oif_aelse_acc_nl;
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl[23:0] = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_10_nl;
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl[23:0] = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_4_nl;
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl[23:0] = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_6_nl;
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl[23:0] = FpAdd_8U_23U_is_a_greater_oif_aelse_acc_8_nl;
  assign nl_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl[7:0] = FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_nl;
  assign nl_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0[7:0] = FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_itm_8_1_mx0w0;
  assign nl_NV_NVDLA_SDP_CORE_Y_idx_core_chn_lut_out_rsci_inst_chn_lut_out_rsci_d = { chn_lut_out_rsci_d_323, chn_lut_out_rsci_d_322, chn_lut_out_rsci_d_321, chn_lut_out_rsci_d_320, chn_lut_out_rsci_d_319, chn_lut_out_rsci_d_318, chn_lut_out_rsci_d_317, chn_lut_out_rsci_d_316, chn_lut_out_rsci_d_315, chn_lut_out_rsci_d_314, chn_lut_out_rsci_d_313, chn_lut_out_rsci_d_312_307, chn_lut_out_rsci_d_306, chn_lut_out_rsci_d_305, chn_lut_out_rsci_d_304, chn_lut_out_rsci_d_303_298, chn_lut_out_rsci_d_297, chn_lut_out_rsci_d_296, chn_lut_out_rsci_d_295, chn_lut_out_rsci_d_294_289, chn_lut_out_rsci_d_288, chn_lut_out_rsci_d_287, chn_lut_out_rsci_d_286, chn_lut_out_rsci_d_285_280, chn_lut_out_rsci_d_279, chn_lut_out_rsci_d_278, chn_lut_out_rsci_d_277, chn_lut_out_rsci_d_276, chn_lut_out_rsci_d_275, chn_lut_out_rsci_d_274, chn_lut_out_rsci_d_273, chn_lut_out_rsci_d_272, chn_lut_out_rsci_d_271, chn_lut_out_rsci_d_270, chn_lut_out_rsci_d_269, chn_lut_out_rsci_d_268, chn_lut_out_rsci_d_267_140, chn_lut_out_rsci_d_139_117, chn_lut_out_rsci_d_116_105, chn_lut_out_rsci_d_104_82, chn_lut_out_rsci_d_81_70, chn_lut_out_rsci_d_69_47, chn_lut_out_rsci_d_46_35, chn_lut_out_rsci_d_34_12, chn_lut_out_rsci_d_11_0 };
  assign nl_acc_10_nl[8:0] = acc_10_nl;
  assign nl_acc_11_nl[8:0] = acc_11_nl;
  assign nl_acc_4_nl[8:0] = acc_4_nl;
  assign nl_acc_5_nl[8:0] = acc_5_nl;
  assign nl_acc_6_nl[8:0] = acc_6_nl;
  assign nl_acc_7_nl[8:0] = acc_7_nl;
  assign nl_acc_8_nl[8:0] = acc_8_nl;
  assign nl_acc_9_nl[8:0] = acc_9_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = { lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, lut_in_data_sva_154[22:0] };
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = { lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] };
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl[49:0] = lut_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl[49:0] = lut_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7:0] = lut_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7:0] = lut_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a = { lut_lookup_1_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2, lut_in_data_sva_154[22:0] };
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl[7:0] = lut_lookup_1_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a = { lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2, cfg_lut_lo_start_1_sva_41[22:0] };
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[4:1] = lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl = lut_lookup_1_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl[49:0] = lut_lookup_1_FpAdd_8U_23U_2_else_2_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl[49:0] = lut_lookup_1_FpAdd_8U_23U_2_if_2_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7:0] = lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl[7:0] = lut_lookup_1_FpAdd_8U_23U_2_if_3_if_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7:0] = lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl[7:0] = lut_lookup_1_FpAdd_8U_23U_2_if_4_if_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = { lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, lut_in_data_sva_154[22:0] };
  assign nl_lut_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = { lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] };
  assign nl_lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1[7:0] = lut_lookup_1_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  assign nl_lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = { lut_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] };
  assign nl_lut_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = { lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] };
  assign nl_lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1[7:0] = lut_lookup_1_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  assign nl_lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl[49:0] = lut_lookup_1_FpAdd_8U_23U_else_2_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl[49:0] = lut_lookup_1_FpAdd_8U_23U_if_2_acc_nl;
  assign nl_lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt[7:0] = lut_lookup_1_FpAdd_8U_23U_if_3_if_acc_sdt;
  assign nl_lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl[7:0] = lut_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a = { 1'b1, FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5 };
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247:0] = lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9:0] = lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a = { 1'b1, FpAdd_8U_23U_2_o_mant_1_lpi_1_dfm_5 };
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a = { 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm };
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247:0] = lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9:0] = lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  assign nl_lut_lookup_1_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a = { 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm };
  assign nl_lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl[22:0] = lut_lookup_1_FpMantRNE_49U_24U_2_else_acc_nl;
  assign nl_lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl[22:0] = lut_lookup_1_FpMantRNE_49U_24U_else_acc_1_nl;
  assign nl_lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl[8:0] = lut_lookup_1_FpNormalize_8U_49U_1_acc_1_nl;
  assign nl_lut_lookup_1_FpNormalize_8U_49U_2_acc_nl[8:0] = lut_lookup_1_FpNormalize_8U_49U_2_acc_nl;
  assign nl_lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl[7:0] = lut_lookup_1_FpNormalize_8U_49U_2_else_acc_nl;
  assign nl_lut_lookup_1_FpNormalize_8U_49U_2_else_lshift_rg_a = FpAdd_8U_23U_2_int_mant_p1_1_sva_3[48:0];
  assign nl_lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt[7:0] = lut_lookup_1_FpNormalize_8U_49U_else_acc_sdt;
  assign nl_lut_lookup_1_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:0];
  assign nl_lut_lookup_1_IntLog2_32U_acc_1_nl[30:0] = lut_lookup_1_IntLog2_32U_acc_1_nl;
  assign nl_lut_lookup_1_IntLog2_32U_lshift_rg_s[31:5] = { reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_10_1_itm[5] };
  assign nl_lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a = { lut_lookup_else_1_lo_index_u_1_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_lut_lookup_1_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a = { lut_lookup_else_else_else_le_index_u_1_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_lut_lookup_1_else_1_acc_nl[32:0] = lut_lookup_1_else_1_acc_nl;
  assign nl_lut_lookup_1_else_1_else_else_acc_nl[8:0] = lut_lookup_1_else_1_else_else_acc_nl;
  assign nl_lut_lookup_1_else_1_else_else_lo_data_f_acc_2[31:0] = lut_lookup_1_else_1_else_else_lo_data_f_acc_2;
  assign nl_lut_lookup_1_else_1_else_else_rshift_rg_s = { reg_lut_lookup_1_else_1_else_else_acc_itm, reg_lut_lookup_1_else_1_else_else_acc_1_itm };
  assign nl_lut_lookup_1_else_else_acc_1_nl[32:0] = lut_lookup_1_else_else_acc_1_nl;
  assign nl_lut_lookup_1_else_else_else_else_acc_itm_mx0w0[8:0] = lut_lookup_1_else_else_else_else_acc_itm_mx0w0;
  assign nl_lut_lookup_1_else_else_else_else_le_data_f_acc_2[31:0] = lut_lookup_1_else_else_else_else_le_data_f_acc_2;
  assign nl_lut_lookup_1_else_else_else_else_rshift_rg_a = { lut_lookup_1_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_1_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_1_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_1_else_else_else_else_le_data_f_and_itm_2 };
  assign nl_lut_lookup_1_else_else_else_else_rshift_rg_s = { reg_lut_lookup_1_else_else_else_else_acc_reg, reg_lut_lookup_1_else_else_else_else_acc_1_reg, reg_lut_lookup_1_else_else_else_else_acc_2_reg, reg_lut_lookup_1_else_else_else_else_acc_3_reg };
  assign nl_lut_lookup_1_else_else_else_if_acc_nl[3:0] = lut_lookup_1_else_else_else_if_acc_nl;
  assign nl_lut_lookup_1_else_if_else_if_acc_nl[3:0] = lut_lookup_1_else_if_else_if_acc_nl;
  assign nl_lut_lookup_1_if_else_else_acc_nl[10:0] = lut_lookup_1_if_else_else_acc_nl;
  assign nl_lut_lookup_1_if_else_else_else_else_acc_nl[32:0] = lut_lookup_1_if_else_else_else_else_acc_nl;
  assign nl_lut_lookup_1_if_else_else_else_else_else_acc_nl[6:0] = lut_lookup_1_if_else_else_else_else_else_acc_nl;
  assign nl_lut_lookup_1_if_else_else_else_else_else_rshift_rg_a = { reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm, reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm };
  assign nl_lut_lookup_1_if_else_else_else_else_else_rshift_rg_s = { reg_lut_lookup_1_else_else_else_else_acc_2_reg, reg_lut_lookup_1_else_else_else_else_acc_3_reg };
  assign nl_lut_lookup_1_if_else_else_else_else_if_acc_nl[3:0] = lut_lookup_1_if_else_else_else_else_if_acc_nl;
  assign nl_lut_lookup_1_if_else_else_else_else_if_lshift_rg_a = { reg_IntLog2_32U_ac_int_cctor_1_30_0_1_itm, reg_IntLog2_32U_ac_int_cctor_1_30_0_1_2_itm };
  assign nl_lut_lookup_1_if_else_else_else_else_if_lshift_rg_s = { reg_lut_lookup_1_else_else_else_else_acc_3_reg, lut_lookup_1_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 };
  assign nl_lut_lookup_1_if_else_else_else_if_acc_nl[3:0] = lut_lookup_1_if_else_else_else_if_acc_nl;
  assign nl_lut_lookup_1_if_if_else_acc_nl[9:0] = lut_lookup_1_if_if_else_acc_nl;
  assign nl_lut_lookup_1_if_if_else_else_if_acc_nl[3:0] = lut_lookup_1_if_if_else_else_if_acc_nl;
  assign nl_lut_lookup_1_leading_sign_49_0_2_rg_mantissa = FpAdd_8U_23U_2_int_mant_p1_1_sva_3[48:0];
  assign nl_lut_lookup_1_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:0];
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = { lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, lut_in_data_sva_154[54:32] };
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = { lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] };
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl[49:0] = lut_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl[49:0] = lut_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7:0] = lut_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7:0] = lut_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a = { lut_lookup_2_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2, lut_in_data_sva_154[54:32] };
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl[7:0] = lut_lookup_2_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a = { lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2, cfg_lut_lo_start_1_sva_41[22:0] };
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl[7:0] = lut_lookup_2_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl[49:0] = lut_lookup_2_FpAdd_8U_23U_2_else_2_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl[49:0] = lut_lookup_2_FpAdd_8U_23U_2_if_2_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7:0] = lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl[7:0] = lut_lookup_2_FpAdd_8U_23U_2_if_3_if_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7:0] = lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl[7:0] = lut_lookup_2_FpAdd_8U_23U_2_if_4_if_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = { lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, lut_in_data_sva_154[54:32] };
  assign nl_lut_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = { lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] };
  assign nl_lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1[7:0] = lut_lookup_2_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  assign nl_lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = { lut_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] };
  assign nl_lut_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = { lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] };
  assign nl_lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1[7:0] = lut_lookup_2_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  assign nl_lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl[49:0] = lut_lookup_2_FpAdd_8U_23U_else_2_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl[49:0] = lut_lookup_2_FpAdd_8U_23U_if_2_acc_nl;
  assign nl_lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt[7:0] = lut_lookup_2_FpAdd_8U_23U_if_3_if_acc_sdt;
  assign nl_lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl[7:0] = lut_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a = { 1'b1, FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5 };
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247:0] = lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9:0] = lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a = { 1'b1, FpAdd_8U_23U_2_o_mant_2_lpi_1_dfm_5 };
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a = { 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg };
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247:0] = lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9:0] = lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  assign nl_lut_lookup_2_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a = { 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg };
  assign nl_lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl[22:0] = lut_lookup_2_FpMantRNE_49U_24U_2_else_acc_nl;
  assign nl_lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl[22:0] = lut_lookup_2_FpMantRNE_49U_24U_else_acc_1_nl;
  assign nl_lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl[8:0] = lut_lookup_2_FpNormalize_8U_49U_1_acc_1_nl;
  assign nl_lut_lookup_2_FpNormalize_8U_49U_2_acc_nl[8:0] = lut_lookup_2_FpNormalize_8U_49U_2_acc_nl;
  assign nl_lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl[7:0] = lut_lookup_2_FpNormalize_8U_49U_2_else_acc_nl;
  assign nl_lut_lookup_2_FpNormalize_8U_49U_2_else_lshift_rg_a = FpAdd_8U_23U_2_int_mant_p1_2_sva_3[48:0];
  assign nl_lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt[7:0] = lut_lookup_2_FpNormalize_8U_49U_else_acc_sdt;
  assign nl_lut_lookup_2_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:0];
  assign nl_lut_lookup_2_IntLog2_32U_acc_1_nl[30:0] = lut_lookup_2_IntLog2_32U_acc_1_nl;
  assign nl_lut_lookup_2_IntLog2_32U_lshift_rg_s[31:5] = { reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_10_1_itm[5] };
  assign nl_lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a = { lut_lookup_else_1_lo_index_u_2_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_lut_lookup_2_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a = { lut_lookup_else_else_else_le_index_u_2_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_lut_lookup_2_else_1_acc_nl[32:0] = lut_lookup_2_else_1_acc_nl;
  assign nl_lut_lookup_2_else_1_else_else_rshift_rg_s = { reg_lut_lookup_2_else_1_else_else_acc_itm, reg_lut_lookup_2_else_1_else_else_acc_1_itm };
  assign nl_lut_lookup_2_else_else_acc_1_nl[32:0] = lut_lookup_2_else_else_acc_1_nl;
  assign nl_lut_lookup_2_else_else_else_else_rshift_rg_a = { lut_lookup_2_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_2_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_2_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_2_else_else_else_else_le_data_f_and_itm_2 };
  assign nl_lut_lookup_2_else_else_else_else_rshift_rg_s = { reg_lut_lookup_2_else_else_else_else_acc_reg, reg_lut_lookup_2_else_else_else_else_acc_1_reg, reg_lut_lookup_2_else_else_else_else_acc_2_reg, reg_lut_lookup_2_else_else_else_else_acc_3_reg };
  assign nl_lut_lookup_2_else_else_else_if_acc_nl[3:0] = lut_lookup_2_else_else_else_if_acc_nl;
  assign nl_lut_lookup_2_else_if_else_if_acc_nl[3:0] = lut_lookup_2_else_if_else_if_acc_nl;
  assign nl_lut_lookup_2_if_else_else_acc_nl[10:0] = lut_lookup_2_if_else_else_acc_nl;
  assign nl_lut_lookup_2_if_else_else_else_else_acc_nl[32:0] = lut_lookup_2_if_else_else_else_else_acc_nl;
  assign nl_lut_lookup_2_if_else_else_else_else_else_acc_nl[6:0] = lut_lookup_2_if_else_else_else_else_else_acc_nl;
  assign nl_lut_lookup_2_if_else_else_else_else_else_rshift_rg_a = { reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg };
  assign nl_lut_lookup_2_if_else_else_else_else_else_rshift_rg_s = { reg_lut_lookup_2_else_else_else_else_acc_2_reg, reg_lut_lookup_2_else_else_else_else_acc_3_reg };
  assign nl_lut_lookup_2_if_else_else_else_else_if_acc_nl[3:0] = lut_lookup_2_if_else_else_else_else_if_acc_nl;
  assign nl_lut_lookup_2_if_else_else_else_else_if_lshift_rg_a = { reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_2_reg };
  assign nl_lut_lookup_2_if_else_else_else_else_if_lshift_rg_s = { reg_lut_lookup_2_else_else_else_else_acc_3_reg, lut_lookup_2_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 };
  assign nl_lut_lookup_2_if_else_else_else_if_acc_nl[3:0] = lut_lookup_2_if_else_else_else_if_acc_nl;
  assign nl_lut_lookup_2_if_if_else_acc_nl[9:0] = lut_lookup_2_if_if_else_acc_nl;
  assign nl_lut_lookup_2_if_if_else_else_if_acc_nl[3:0] = lut_lookup_2_if_if_else_else_if_acc_nl;
  assign nl_lut_lookup_2_leading_sign_49_0_2_rg_mantissa = FpAdd_8U_23U_2_int_mant_p1_2_sva_3[48:0];
  assign nl_lut_lookup_2_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:0];
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = { lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, lut_in_data_sva_154[86:64] };
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = { lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] };
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl[49:0] = lut_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl[49:0] = lut_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7:0] = lut_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7:0] = lut_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a = { lut_lookup_3_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2, lut_in_data_sva_154[86:64] };
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl[7:0] = lut_lookup_3_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a = { lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2, cfg_lut_lo_start_1_sva_41[22:0] };
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl[7:0] = lut_lookup_3_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl[49:0] = lut_lookup_3_FpAdd_8U_23U_2_else_2_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl[49:0] = lut_lookup_3_FpAdd_8U_23U_2_if_2_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7:0] = lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl[7:0] = lut_lookup_3_FpAdd_8U_23U_2_if_3_if_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7:0] = lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl[7:0] = lut_lookup_3_FpAdd_8U_23U_2_if_4_if_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = { lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, lut_in_data_sva_154[86:64] };
  assign nl_lut_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = { lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] };
  assign nl_lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1[7:0] = lut_lookup_3_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  assign nl_lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = { lut_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] };
  assign nl_lut_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = { lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] };
  assign nl_lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1[7:0] = lut_lookup_3_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  assign nl_lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl[49:0] = lut_lookup_3_FpAdd_8U_23U_else_2_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl[49:0] = lut_lookup_3_FpAdd_8U_23U_if_2_acc_nl;
  assign nl_lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt[7:0] = lut_lookup_3_FpAdd_8U_23U_if_3_if_acc_sdt;
  assign nl_lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl[7:0] = lut_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a = { 1'b1, FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5 };
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247:0] = lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9:0] = lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a = { 1'b1, FpAdd_8U_23U_2_o_mant_3_lpi_1_dfm_5 };
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a = { 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg };
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247:0] = lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9:0] = lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  assign nl_lut_lookup_3_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a = { 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg };
  assign nl_lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl[22:0] = lut_lookup_3_FpMantRNE_49U_24U_2_else_acc_nl;
  assign nl_lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl[22:0] = lut_lookup_3_FpMantRNE_49U_24U_else_acc_1_nl;
  assign nl_lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl[8:0] = lut_lookup_3_FpNormalize_8U_49U_1_acc_1_nl;
  assign nl_lut_lookup_3_FpNormalize_8U_49U_2_acc_nl[8:0] = lut_lookup_3_FpNormalize_8U_49U_2_acc_nl;
  assign nl_lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl[7:0] = lut_lookup_3_FpNormalize_8U_49U_2_else_acc_nl;
  assign nl_lut_lookup_3_FpNormalize_8U_49U_2_else_lshift_rg_a = FpAdd_8U_23U_2_int_mant_p1_3_sva_3[48:0];
  assign nl_lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt[7:0] = lut_lookup_3_FpNormalize_8U_49U_else_acc_sdt;
  assign nl_lut_lookup_3_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:0];
  assign nl_lut_lookup_3_IntLog2_32U_acc_1_nl[30:0] = lut_lookup_3_IntLog2_32U_acc_1_nl;
  assign nl_lut_lookup_3_IntLog2_32U_lshift_rg_s[31:5] = { reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_10_1_itm[5] };
  assign nl_lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a = { lut_lookup_else_1_lo_index_u_3_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_lut_lookup_3_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a = { lut_lookup_else_else_else_le_index_u_3_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_lut_lookup_3_else_1_acc_nl[32:0] = lut_lookup_3_else_1_acc_nl;
  assign nl_lut_lookup_3_else_1_else_else_rshift_rg_s = { reg_lut_lookup_3_else_1_else_else_acc_itm, reg_lut_lookup_3_else_1_else_else_acc_1_itm };
  assign nl_lut_lookup_3_else_else_acc_1_nl[32:0] = lut_lookup_3_else_else_acc_1_nl;
  assign nl_lut_lookup_3_else_else_else_else_rshift_rg_a = { lut_lookup_3_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_3_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_3_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_3_else_else_else_else_le_data_f_and_itm_2 };
  assign nl_lut_lookup_3_else_else_else_else_rshift_rg_s = { reg_lut_lookup_3_else_else_else_else_acc_reg, reg_lut_lookup_3_else_else_else_else_acc_1_reg, reg_lut_lookup_3_else_else_else_else_acc_2_reg, reg_lut_lookup_3_else_else_else_else_acc_3_reg };
  assign nl_lut_lookup_3_else_else_else_if_acc_nl[3:0] = lut_lookup_3_else_else_else_if_acc_nl;
  assign nl_lut_lookup_3_else_if_else_if_acc_nl[3:0] = lut_lookup_3_else_if_else_if_acc_nl;
  assign nl_lut_lookup_3_if_else_else_acc_nl[10:0] = lut_lookup_3_if_else_else_acc_nl;
  assign nl_lut_lookup_3_if_else_else_else_else_acc_nl[32:0] = lut_lookup_3_if_else_else_else_else_acc_nl;
  assign nl_lut_lookup_3_if_else_else_else_else_else_acc_nl[6:0] = lut_lookup_3_if_else_else_else_else_else_acc_nl;
  assign nl_lut_lookup_3_if_else_else_else_else_else_rshift_rg_a = { reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg };
  assign nl_lut_lookup_3_if_else_else_else_else_else_rshift_rg_s = { reg_lut_lookup_3_else_else_else_else_acc_2_reg, reg_lut_lookup_3_else_else_else_else_acc_3_reg };
  assign nl_lut_lookup_3_if_else_else_else_else_if_acc_nl[3:0] = lut_lookup_3_if_else_else_else_else_if_acc_nl;
  assign nl_lut_lookup_3_if_else_else_else_else_if_lshift_rg_a = { reg_IntLog2_32U_ac_int_cctor_1_30_0_3_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_3_2_reg };
  assign nl_lut_lookup_3_if_else_else_else_else_if_lshift_rg_s = { reg_lut_lookup_3_else_else_else_else_acc_3_reg, lut_lookup_3_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 };
  assign nl_lut_lookup_3_if_else_else_else_if_acc_nl[3:0] = lut_lookup_3_if_else_else_else_if_acc_nl;
  assign nl_lut_lookup_3_if_if_else_acc_nl[9:0] = lut_lookup_3_if_if_else_acc_nl;
  assign nl_lut_lookup_3_if_if_else_else_if_acc_nl[3:0] = lut_lookup_3_if_if_else_else_if_acc_nl;
  assign nl_lut_lookup_3_leading_sign_49_0_2_rg_mantissa = FpAdd_8U_23U_2_int_mant_p1_3_sva_3[48:0];
  assign nl_lut_lookup_3_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:0];
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = { lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, lut_in_data_sva_154[118:96] };
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = { lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] };
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl[49:0] = lut_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl[49:0] = lut_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl[7:0] = lut_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_2_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl[7:0] = lut_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_2_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_a = { lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_6_or_itm_2, lut_in_data_sva_154[118:96] };
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_a_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl[7:0] = lut_lookup_4_FpAdd_8U_23U_2_a_left_shift_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_a = { lut_lookup_4_FpAdd_8U_23U_2_IsZero_8U_23U_7_or_itm_2, cfg_lut_lo_start_1_sva_41[22:0] };
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_b_int_mant_p1_lshift_rg_s[8:1] = lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl[7:0] = lut_lookup_4_FpAdd_8U_23U_2_b_left_shift_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl[49:0] = lut_lookup_4_FpAdd_8U_23U_2_else_2_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl[49:0] = lut_lookup_4_FpAdd_8U_23U_2_if_2_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl[7:0] = lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_1_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl[7:0] = lut_lookup_4_FpAdd_8U_23U_2_if_3_if_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl[7:0] = lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_1_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl[7:0] = lut_lookup_4_FpAdd_8U_23U_2_if_4_if_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = { lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_4_or_itm_2, lut_in_data_sva_154[118:96] };
  assign nl_lut_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = { lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1, nl_lut_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[0] };
  assign nl_lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1[7:0] = lut_lookup_4_FpAdd_8U_23U_a_left_shift_conc_6_8_1;
  assign nl_lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = { lut_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2, cfg_lut_le_start_1_sva_41[22:0] };
  assign nl_lut_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = { lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1, nl_lut_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[0] };
  assign nl_lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1[7:0] = lut_lookup_4_FpAdd_8U_23U_b_left_shift_conc_6_8_1;
  assign nl_lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl[49:0] = lut_lookup_4_FpAdd_8U_23U_else_2_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl[49:0] = lut_lookup_4_FpAdd_8U_23U_if_2_acc_nl;
  assign nl_lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt[7:0] = lut_lookup_4_FpAdd_8U_23U_if_3_if_acc_sdt;
  assign nl_lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl[7:0] = lut_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_else_lshift_rg_a = { 1'b1, FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5 };
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl[247:0] = lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_if_1_acc_nl;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp[9:0] = lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_lshift_acc_tmp;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_1_m_int_lshift_rg_a = { 1'b1, FpAdd_8U_23U_2_o_mant_lpi_1_dfm_5 };
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_else_lshift_rg_a = { 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 };
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl[247:0] = lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_if_1_acc_nl;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp[9:0] = lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_lshift_acc_tmp;
  assign nl_lut_lookup_4_FpFloatToIntFrac_8U_23U_8U_9U_35U_m_int_lshift_rg_a = { 1'b1, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 };
  assign nl_lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl[22:0] = lut_lookup_4_FpMantRNE_49U_24U_2_else_acc_nl;
  assign nl_lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl[22:0] = lut_lookup_4_FpMantRNE_49U_24U_else_acc_1_nl;
  assign nl_lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl[8:0] = lut_lookup_4_FpNormalize_8U_49U_1_acc_1_nl;
  assign nl_lut_lookup_4_FpNormalize_8U_49U_2_acc_nl[8:0] = lut_lookup_4_FpNormalize_8U_49U_2_acc_nl;
  assign nl_lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl[7:0] = lut_lookup_4_FpNormalize_8U_49U_2_else_acc_nl;
  assign nl_lut_lookup_4_FpNormalize_8U_49U_2_else_lshift_rg_a = FpAdd_8U_23U_2_int_mant_p1_sva_3[48:0];
  assign nl_lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt[7:0] = lut_lookup_4_FpNormalize_8U_49U_else_acc_sdt;
  assign nl_lut_lookup_4_FpNormalize_8U_49U_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_sva_3[48:0];
  assign nl_lut_lookup_4_IntLog2_32U_acc_1_nl[30:0] = lut_lookup_4_IntLog2_32U_acc_1_nl;
  assign nl_lut_lookup_4_IntLog2_32U_lshift_rg_s[31:5] = { reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5], reg_FpAdd_8U_23U_1_o_expo_lpi_1_dfm_10_1_itm[5] };
  assign nl_lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_1_mbits_fixed_rshift_rg_a = { lut_lookup_else_1_lo_index_u_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_lut_lookup_4_IntSignedShiftRightTZ_32U_8U_9U_mbits_fixed_rshift_rg_a = { lut_lookup_else_else_else_le_index_u_sva_3, 127'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 };
  assign nl_lut_lookup_4_else_1_acc_nl[32:0] = lut_lookup_4_else_1_acc_nl;
  assign nl_lut_lookup_4_else_1_else_else_rshift_rg_s = { reg_lut_lookup_4_else_1_else_else_acc_itm, reg_lut_lookup_4_else_1_else_else_acc_1_itm };
  assign nl_lut_lookup_4_else_else_acc_1_nl[32:0] = lut_lookup_4_else_else_acc_1_nl;
  assign nl_lut_lookup_4_else_else_else_else_rshift_rg_a = { lut_lookup_4_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_4_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_4_else_else_else_else_le_data_f_and_itm_2[31], lut_lookup_4_else_else_else_else_le_data_f_and_itm_2 };
  assign nl_lut_lookup_4_else_else_else_else_rshift_rg_s = { reg_lut_lookup_4_else_else_else_else_acc_reg, reg_lut_lookup_4_else_else_else_else_acc_1_reg, reg_lut_lookup_4_else_else_else_else_acc_2_reg, reg_lut_lookup_4_else_else_else_else_acc_3_reg };
  assign nl_lut_lookup_4_else_else_else_if_acc_nl[3:0] = lut_lookup_4_else_else_else_if_acc_nl;
  assign nl_lut_lookup_4_else_if_else_if_acc_nl[3:0] = lut_lookup_4_else_if_else_if_acc_nl;
  assign nl_lut_lookup_4_if_else_else_acc_nl[10:0] = lut_lookup_4_if_else_else_acc_nl;
  assign nl_lut_lookup_4_if_else_else_else_else_acc_nl[32:0] = lut_lookup_4_if_else_else_else_else_acc_nl;
  assign nl_lut_lookup_4_if_else_else_else_else_else_acc_nl[6:0] = lut_lookup_4_if_else_else_else_else_else_acc_nl;
  assign nl_lut_lookup_4_if_else_else_else_else_else_rshift_rg_a = { reg_IntLog2_32U_ac_int_cctor_1_30_0_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 };
  assign nl_lut_lookup_4_if_else_else_else_else_else_rshift_rg_s = { reg_lut_lookup_4_else_else_else_else_acc_2_reg, reg_lut_lookup_4_else_else_else_else_acc_3_reg };
  assign nl_lut_lookup_4_if_else_else_else_else_if_acc_nl[3:0] = lut_lookup_4_if_else_else_else_else_if_acc_nl;
  assign nl_lut_lookup_4_if_else_else_else_else_if_lshift_rg_a = { reg_IntLog2_32U_ac_int_cctor_1_30_0_reg, reg_IntLog2_32U_ac_int_cctor_1_30_0_2_reg_1 };
  assign nl_lut_lookup_4_if_else_else_else_else_if_lshift_rg_s = { reg_lut_lookup_4_else_else_else_else_acc_3_reg, lut_lookup_4_IntLog2_32U_leadzero_slc_IntLog2_32U_leadzero_5_0_4_0_6_itm_3 };
  assign nl_lut_lookup_4_if_else_else_else_if_acc_nl[3:0] = lut_lookup_4_if_else_else_else_if_acc_nl;
  assign nl_lut_lookup_4_if_if_else_acc_nl[9:0] = lut_lookup_4_if_if_else_acc_nl;
  assign nl_lut_lookup_4_if_if_else_else_if_acc_nl[3:0] = lut_lookup_4_if_if_else_else_if_acc_nl;
  assign nl_lut_lookup_4_leading_sign_49_0_2_rg_mantissa = FpAdd_8U_23U_2_int_mant_p1_sva_3[48:0];
  assign nl_lut_lookup_4_leading_sign_49_0_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_sva_3[48:0];
  assign nl_lut_lookup_if_else_else_else_le_index_s_1_sva[8:0] = lut_lookup_if_else_else_else_le_index_s_1_sva;
  assign nl_lut_lookup_if_else_else_else_le_index_s_2_sva[8:0] = lut_lookup_if_else_else_else_le_index_s_2_sva;
  assign nl_lut_lookup_if_else_else_else_le_index_s_3_sva[8:0] = lut_lookup_if_else_else_else_le_index_s_3_sva;
  assign nl_lut_lookup_if_else_else_else_le_index_s_sva[8:0] = lut_lookup_if_else_else_else_le_index_s_sva;
  assign nl_lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0[31:0] = lut_lookup_if_else_else_le_data_sub_1_sva_mx0w0;
  assign nl_lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0[31:0] = lut_lookup_if_else_else_le_data_sub_2_sva_mx0w0;
  assign nl_lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0[31:0] = lut_lookup_if_else_else_le_data_sub_3_sva_mx0w0;
  assign nl_lut_lookup_if_else_else_le_data_sub_sva_mx0w0[31:0] = lut_lookup_if_else_else_le_data_sub_sva_mx0w0;
  assign nl_lut_lookup_if_if_else_else_le_index_s_1_sva[8:0] = lut_lookup_if_if_else_else_le_index_s_1_sva;
  assign nl_lut_lookup_if_if_else_else_le_index_s_2_sva[8:0] = lut_lookup_if_if_else_else_le_index_s_2_sva;
  assign nl_lut_lookup_if_if_else_else_le_index_s_3_sva[8:0] = lut_lookup_if_if_else_else_le_index_s_3_sva;
  assign nl_lut_lookup_if_if_else_else_le_index_s_sva[8:0] = lut_lookup_if_if_else_else_le_index_s_sva;
  assign nl_z_out_4[8:0] = z_out_4;
  assign nl_z_out_5[8:0] = z_out_5;
  assign nl_z_out_6[8:0] = z_out_6;
  assign nl_z_out_7[8:0] = z_out_7;
  assign or_1691_cse = or_1688_cse;
endmodule
