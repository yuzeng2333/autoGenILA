module \$paramod\SDP_Y_CORE_mgc_in_wire_v1\rscid=18\width=2 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:376" *)
  output [1:0] d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:377" *)
  input [1:0] z;
  assign d = z;
endmodule
