module \$paramod\SDP_Y_CORE_mgc_in_wire_v1\rscid=4\width=1 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:376" *)
  output d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_core.v:377" *)
  input z;
  assign d = z;
endmodule
