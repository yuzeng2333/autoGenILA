module aes_s(clk, in, out);
  wire [7:0] _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  input clk;
  input [7:0] in;
  output [7:0] out;
  reg [7:0] out;
  always @(posedge clk)
      out <= _000_;
  assign _001_ = in == 8'h9e;
  assign _002_ = in == 8'h9d;
  assign _003_ = in == 8'h9c;
  assign _004_ = in == 8'h9b;
  assign _005_ = in == 8'h9a;
  assign _006_ = in == 8'h99;
  assign _007_ = in == 8'h98;
  assign _008_ = in == 8'h97;
  assign _009_ = in == 8'h96;
  assign _010_ = in == 8'h95;
  assign _011_ = in == 8'hf8;
  assign _012_ = in == 8'h94;
  assign _013_ = in == 8'h93;
  assign _014_ = in == 8'h92;
  assign _015_ = in == 8'h91;
  assign _016_ = in == 8'h90;
  assign _017_ = in == 8'h8f;
  assign _018_ = in == 8'h8e;
  assign _019_ = in == 8'h8d;
  assign _020_ = in == 8'h8c;
  assign _021_ = in == 8'h8b;
  assign _022_ = in == 8'hf7;
  assign _023_ = in == 8'h8a;
  assign _024_ = in == 8'h89;
  assign _025_ = in == 8'h88;
  assign _026_ = in == 8'h87;
  assign _027_ = in == 8'h86;
  assign _028_ = in == 8'h85;
  assign _029_ = in == 8'h84;
  assign _030_ = in == 8'h83;
  assign _031_ = in == 8'h82;
  assign _032_ = in == 8'h81;
  assign _033_ = in == 8'hf6;
  assign _034_ = in == 8'h80;
  assign _035_ = in == 7'h7f;
  assign _036_ = in == 7'h7e;
  assign _037_ = in == 7'h7d;
  assign _038_ = in == 7'h7c;
  assign _039_ = in == 7'h7b;
  assign _040_ = in == 7'h7a;
  assign _041_ = in == 7'h79;
  assign _042_ = in == 7'h78;
  assign _043_ = in == 7'h77;
  assign _044_ = in == 8'hf5;
  assign _045_ = in == 7'h76;
  assign _046_ = in == 7'h75;
  assign _047_ = in == 7'h74;
  assign _048_ = in == 7'h73;
  assign _049_ = in == 7'h72;
  assign _050_ = in == 7'h71;
  assign _051_ = in == 7'h70;
  assign _052_ = in == 7'h6f;
  assign _053_ = in == 7'h6e;
  assign _054_ = in == 7'h6d;
  assign _055_ = in == 8'hf4;
  assign _056_ = in == 7'h6c;
  assign _057_ = in == 7'h6b;
  assign _058_ = in == 7'h6a;
  assign _059_ = in == 7'h69;
  assign _060_ = in == 7'h68;
  assign _061_ = in == 7'h67;
  assign _062_ = in == 7'h66;
  assign _063_ = in == 7'h65;
  assign _064_ = in == 7'h64;
  assign _065_ = in == 7'h63;
  assign _066_ = in == 8'hf3;
  assign _067_ = in == 7'h62;
  assign _068_ = in == 7'h61;
  assign _069_ = in == 7'h60;
  assign _070_ = in == 7'h5f;
  assign _071_ = in == 7'h5e;
  assign _072_ = in == 7'h5d;
  assign _073_ = in == 7'h5c;
  assign _074_ = in == 7'h5b;
  assign _075_ = in == 7'h5a;
  assign _076_ = in == 7'h59;
  assign _077_ = in == 8'hf2;
  assign _078_ = in == 7'h58;
  assign _079_ = in == 7'h57;
  assign _080_ = in == 7'h56;
  assign _081_ = in == 7'h55;
  assign _082_ = in == 7'h54;
  assign _083_ = in == 7'h53;
  assign _084_ = in == 7'h52;
  assign _085_ = in == 7'h51;
  assign _086_ = in == 7'h50;
  assign _087_ = in == 7'h4f;
  assign _088_ = in == 8'hf1;
  assign _089_ = in == 7'h4e;
  assign _090_ = in == 7'h4d;
  assign _091_ = in == 7'h4c;
  assign _092_ = in == 7'h4b;
  assign _093_ = in == 7'h4a;
  assign _094_ = in == 7'h49;
  assign _095_ = in == 7'h48;
  assign _096_ = in == 7'h47;
  assign _097_ = in == 7'h46;
  assign _098_ = in == 7'h45;
  assign _099_ = in == 8'hf0;
  assign _100_ = in == 7'h44;
  assign _101_ = in == 7'h43;
  assign _102_ = in == 7'h42;
  assign _103_ = in == 7'h41;
  assign _104_ = in == 7'h40;
  assign _105_ = in == 6'h3f;
  assign _106_ = in == 6'h3e;
  assign _107_ = in == 6'h3d;
  assign _108_ = in == 6'h3c;
  assign _109_ = in == 6'h3b;
  assign _110_ = in == 8'hef;
  wire [255:0] fangyuan0;
  assign fangyuan0 = { _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_, _156_, _155_, _153_, _152_, _151_, _150_, _149_, _148_, _147_, _146_, _145_, _144_, _142_, _141_, _140_, _139_, _138_, _137_, _136_, _135_, _134_, _133_, _131_, _130_, _129_, _128_, _127_, _126_, _125_, _124_, _123_, _122_, _120_, _119_, _118_, _117_, _116_, _115_, _114_, _113_, _112_, _111_, _109_, _108_, _107_, _106_, _105_, _104_, _103_, _102_, _101_, _100_, _098_, _097_, _096_, _095_, _094_, _093_, _092_, _091_, _090_, _089_, _087_, _086_, _085_, _084_, _083_, _082_, _081_, _080_, _079_, _078_, _076_, _075_, _074_, _073_, _072_, _071_, _070_, _069_, _068_, _067_, _065_, _064_, _063_, _062_, _061_, _060_, _059_, _058_, _057_, _056_, _054_, _053_, _052_, _051_, _050_, _049_, _048_, _047_, _046_, _045_, _043_, _042_, _041_, _040_, _039_, _038_, _037_, _036_, _035_, _034_, _032_, _031_, _030_, _029_, _028_, _027_, _026_, _025_, _024_, _023_, _021_, _020_, _019_, _018_, _017_, _016_, _015_, _014_, _013_, _012_, _010_, _009_, _008_, _007_, _006_, _005_, _004_, _003_, _002_, _001_, _255_, _254_, _253_, _252_, _251_, _250_, _249_, _248_, _247_, _246_, _244_, _243_, _242_, _241_, _240_, _239_, _238_, _237_, _236_, _235_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_, _214_, _213_, _211_, _210_, _209_, _208_, _207_, _206_, _205_, _204_, _203_, _202_, _200_, _199_, _198_, _197_, _196_, _195_, _194_, _193_, _192_, _191_, _189_, _188_, _187_, _186_, _185_, _184_, _183_, _182_, _181_, _180_, _179_, _178_, _177_, _176_, _175_, _165_, _154_, _143_, _132_, _121_, _110_, _099_, _088_, _077_, _066_, _055_, _044_, _033_, _022_, _011_, _256_, _245_, _234_, _223_, _212_, _201_, _190_ };

  always @(out or fangyuan0) begin
    casez (fangyuan0)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _000_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _000_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _000_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _000_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _000_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _000_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _000_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _000_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _000_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _000_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _000_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _000_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _000_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _000_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _000_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _000_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _000_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _000_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _000_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _000_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _000_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _000_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _000_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _000_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _000_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _000_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _000_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _000_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _000_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _000_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _000_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _000_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _000_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _000_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _000_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _000_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _000_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _000_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _000_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _000_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _000_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _000_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _000_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _000_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _000_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _000_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _000_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _000_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _000_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _000_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _000_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _000_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _000_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _000_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _000_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _000_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _000_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _000_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _000_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _000_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _000_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _000_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _000_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100011 ;
      default:
        _000_ = out ;
    endcase
  end
  assign _111_ = in == 6'h3a;
  assign _112_ = in == 6'h39;
  assign _113_ = in == 6'h38;
  assign _114_ = in == 6'h37;
  assign _115_ = in == 6'h36;
  assign _116_ = in == 6'h35;
  assign _117_ = in == 6'h34;
  assign _118_ = in == 6'h33;
  assign _119_ = in == 6'h32;
  assign _120_ = in == 6'h31;
  assign _121_ = in == 8'hee;
  assign _122_ = in == 6'h30;
  assign _123_ = in == 6'h2f;
  assign _124_ = in == 6'h2e;
  assign _125_ = in == 6'h2d;
  assign _126_ = in == 6'h2c;
  assign _127_ = in == 6'h2b;
  assign _128_ = in == 6'h2a;
  assign _129_ = in == 6'h29;
  assign _130_ = in == 6'h28;
  assign _131_ = in == 6'h27;
  assign _132_ = in == 8'hed;
  assign _133_ = in == 6'h26;
  assign _134_ = in == 6'h25;
  assign _135_ = in == 6'h24;
  assign _136_ = in == 6'h23;
  assign _137_ = in == 6'h22;
  assign _138_ = in == 6'h21;
  assign _139_ = in == 6'h20;
  assign _140_ = in == 5'h1f;
  assign _141_ = in == 5'h1e;
  assign _142_ = in == 5'h1d;
  assign _143_ = in == 8'hec;
  assign _144_ = in == 5'h1c;
  assign _145_ = in == 5'h1b;
  assign _146_ = in == 5'h1a;
  assign _147_ = in == 5'h19;
  assign _148_ = in == 5'h18;
  assign _149_ = in == 5'h17;
  assign _150_ = in == 5'h16;
  assign _151_ = in == 5'h15;
  assign _152_ = in == 5'h14;
  assign _153_ = in == 5'h13;
  assign _154_ = in == 8'heb;
  assign _155_ = in == 5'h12;
  assign _156_ = in == 5'h11;
  assign _157_ = in == 5'h10;
  assign _158_ = in == 4'hf;
  assign _159_ = in == 4'he;
  assign _160_ = in == 4'hd;
  assign _161_ = in == 4'hc;
  assign _162_ = in == 4'hb;
  assign _163_ = in == 4'ha;
  assign _164_ = in == 4'h9;
  assign _165_ = in == 8'hea;
  assign _166_ = in == 4'h8;
  assign _167_ = in == 3'h7;
  assign _168_ = in == 3'h6;
  assign _169_ = in == 3'h5;
  assign _170_ = in == 3'h4;
  assign _171_ = in == 2'h3;
  assign _172_ = in == 2'h2;
  assign _173_ = in == 1'h1;
  assign _174_ = ! in;
  assign _175_ = in == 8'he9;
  assign _176_ = in == 8'he8;
  assign _177_ = in == 8'he7;
  assign _178_ = in == 8'he6;
  assign _179_ = in == 8'he5;
  assign _180_ = in == 8'he4;
  assign _181_ = in == 8'he3;
  assign _182_ = in == 8'he2;
  assign _183_ = in == 8'he1;
  assign _184_ = in == 8'he0;
  assign _185_ = in == 8'hdf;
  assign _186_ = in == 8'hde;
  assign _187_ = in == 8'hdd;
  assign _188_ = in == 8'hdc;
  assign _189_ = in == 8'hdb;
  assign _190_ = in == 8'hff;
  assign _191_ = in == 8'hda;
  assign _192_ = in == 8'hd9;
  assign _193_ = in == 8'hd8;
  assign _194_ = in == 8'hd7;
  assign _195_ = in == 8'hd6;
  assign _196_ = in == 8'hd5;
  assign _197_ = in == 8'hd4;
  assign _198_ = in == 8'hd3;
  assign _199_ = in == 8'hd2;
  assign _200_ = in == 8'hd1;
  assign _201_ = in == 8'hfe;
  assign _202_ = in == 8'hd0;
  assign _203_ = in == 8'hcf;
  assign _204_ = in == 8'hce;
  assign _205_ = in == 8'hcd;
  assign _206_ = in == 8'hcc;
  assign _207_ = in == 8'hcb;
  assign _208_ = in == 8'hca;
  assign _209_ = in == 8'hc9;
  assign _210_ = in == 8'hc8;
  assign _211_ = in == 8'hc7;
  assign _212_ = in == 8'hfd;
  assign _213_ = in == 8'hc6;
  assign _214_ = in == 8'hc5;
  assign _215_ = in == 8'hc4;
  assign _216_ = in == 8'hc3;
  assign _217_ = in == 8'hc2;
  assign _218_ = in == 8'hc1;
  assign _219_ = in == 8'hc0;
  assign _220_ = in == 8'hbf;
  assign _221_ = in == 8'hbe;
  assign _222_ = in == 8'hbd;
  assign _223_ = in == 8'hfc;
  assign _224_ = in == 8'hbc;
  assign _225_ = in == 8'hbb;
  assign _226_ = in == 8'hba;
  assign _227_ = in == 8'hb9;
  assign _228_ = in == 8'hb8;
  assign _229_ = in == 8'hb7;
  assign _230_ = in == 8'hb6;
  assign _231_ = in == 8'hb5;
  assign _232_ = in == 8'hb4;
  assign _233_ = in == 8'hb3;
  assign _234_ = in == 8'hfb;
  assign _235_ = in == 8'hb2;
  assign _236_ = in == 8'hb1;
  assign _237_ = in == 8'hb0;
  assign _238_ = in == 8'haf;
  assign _239_ = in == 8'hae;
  assign _240_ = in == 8'had;
  assign _241_ = in == 8'hac;
  assign _242_ = in == 8'hab;
  assign _243_ = in == 8'haa;
  assign _244_ = in == 8'ha9;
  assign _245_ = in == 8'hfa;
  assign _246_ = in == 8'ha8;
  assign _247_ = in == 8'ha7;
  assign _248_ = in == 8'ha6;
  assign _249_ = in == 8'ha5;
  assign _250_ = in == 8'ha4;
  assign _251_ = in == 8'ha3;
  assign _252_ = in == 8'ha2;
  assign _253_ = in == 8'ha1;
  assign _254_ = in == 8'ha0;
  assign _255_ = in == 8'h9f;
  assign _256_ = in == 8'hf9;
endmodule
