module AesDecrypt(clock, reset, io_dataIn, io_ivIn, io_dataValid, io_keys_0_0_0, io_keys_0_0_1, io_keys_0_0_2, io_keys_0_0_3, io_keys_0_1_0, io_keys_0_1_1, io_keys_0_1_2, io_keys_0_1_3, io_keys_0_2_0, io_keys_0_2_1, io_keys_0_2_2, io_keys_0_2_3, io_keys_0_3_0, io_keys_0_3_1, io_keys_0_3_2, io_keys_0_3_3, io_keys_1_0_0, io_keys_1_0_1, io_keys_1_0_2, io_keys_1_0_3, io_keys_1_1_0, io_keys_1_1_1, io_keys_1_1_2, io_keys_1_1_3, io_keys_1_2_0, io_keys_1_2_1, io_keys_1_2_2, io_keys_1_2_3, io_keys_1_3_0, io_keys_1_3_1, io_keys_1_3_2, io_keys_1_3_3, io_keys_2_0_0, io_keys_2_0_1, io_keys_2_0_2, io_keys_2_0_3, io_keys_2_1_0, io_keys_2_1_1, io_keys_2_1_2, io_keys_2_1_3, io_keys_2_2_0, io_keys_2_2_1, io_keys_2_2_2, io_keys_2_2_3, io_keys_2_3_0, io_keys_2_3_1, io_keys_2_3_2, io_keys_2_3_3, io_keys_3_0_0, io_keys_3_0_1, io_keys_3_0_2, io_keys_3_0_3, io_keys_3_1_0, io_keys_3_1_1, io_keys_3_1_2, io_keys_3_1_3, io_keys_3_2_0, io_keys_3_2_1, io_keys_3_2_2, io_keys_3_2_3, io_keys_3_3_0, io_keys_3_3_1, io_keys_3_3_2, io_keys_3_3_3, io_keys_4_0_0, io_keys_4_0_1, io_keys_4_0_2, io_keys_4_0_3, io_keys_4_1_0, io_keys_4_1_1, io_keys_4_1_2, io_keys_4_1_3, io_keys_4_2_0, io_keys_4_2_1, io_keys_4_2_2, io_keys_4_2_3, io_keys_4_3_0, io_keys_4_3_1, io_keys_4_3_2, io_keys_4_3_3, io_keys_5_0_0, io_keys_5_0_1, io_keys_5_0_2, io_keys_5_0_3, io_keys_5_1_0, io_keys_5_1_1, io_keys_5_1_2, io_keys_5_1_3, io_keys_5_2_0, io_keys_5_2_1, io_keys_5_2_2, io_keys_5_2_3, io_keys_5_3_0, io_keys_5_3_1, io_keys_5_3_2, io_keys_5_3_3, io_keys_6_0_0, io_keys_6_0_1, io_keys_6_0_2, io_keys_6_0_3, io_keys_6_1_0, io_keys_6_1_1, io_keys_6_1_2, io_keys_6_1_3, io_keys_6_2_0, io_keys_6_2_1, io_keys_6_2_2, io_keys_6_2_3, io_keys_6_3_0, io_keys_6_3_1, io_keys_6_3_2, io_keys_6_3_3, io_keys_7_0_0, io_keys_7_0_1, io_keys_7_0_2, io_keys_7_0_3, io_keys_7_1_0, io_keys_7_1_1, io_keys_7_1_2, io_keys_7_1_3, io_keys_7_2_0, io_keys_7_2_1, io_keys_7_2_2, io_keys_7_2_3, io_keys_7_3_0, io_keys_7_3_1, io_keys_7_3_2, io_keys_7_3_3, io_keys_8_0_0, io_keys_8_0_1, io_keys_8_0_2, io_keys_8_0_3, io_keys_8_1_0, io_keys_8_1_1, io_keys_8_1_2, io_keys_8_1_3, io_keys_8_2_0, io_keys_8_2_1, io_keys_8_2_2, io_keys_8_2_3, io_keys_8_3_0, io_keys_8_3_1, io_keys_8_3_2, io_keys_8_3_3, io_keys_9_0_0, io_keys_9_0_1, io_keys_9_0_2, io_keys_9_0_3, io_keys_9_1_0, io_keys_9_1_1, io_keys_9_1_2, io_keys_9_1_3, io_keys_9_2_0, io_keys_9_2_1, io_keys_9_2_2, io_keys_9_2_3, io_keys_9_3_0, io_keys_9_3_1, io_keys_9_3_2, io_keys_9_3_3, io_keys_10_0_0, io_keys_10_0_1, io_keys_10_0_2, io_keys_10_0_3, io_keys_10_1_0, io_keys_10_1_1, io_keys_10_1_2, io_keys_10_1_3, io_keys_10_2_0, io_keys_10_2_1, io_keys_10_2_2, io_keys_10_2_3, io_keys_10_3_0, io_keys_10_3_1, io_keys_10_3_2, io_keys_10_3_3, io_keys_11_0_0, io_keys_11_0_1, io_keys_11_0_2, io_keys_11_0_3, io_keys_11_1_0, io_keys_11_1_1, io_keys_11_1_2, io_keys_11_1_3, io_keys_11_2_0, io_keys_11_2_1, io_keys_11_2_2, io_keys_11_2_3, io_keys_11_3_0, io_keys_11_3_1, io_keys_11_3_2, io_keys_11_3_3, io_keys_12_0_0, io_keys_12_0_1, io_keys_12_0_2, io_keys_12_0_3, io_keys_12_1_0, io_keys_12_1_1, io_keys_12_1_2, io_keys_12_1_3, io_keys_12_2_0, io_keys_12_2_1, io_keys_12_2_2, io_keys_12_2_3, io_keys_12_3_0, io_keys_12_3_1, io_keys_12_3_2, io_keys_12_3_3, io_keys_13_0_0, io_keys_13_0_1, io_keys_13_0_2, io_keys_13_0_3, io_keys_13_1_0, io_keys_13_1_1, io_keys_13_1_2, io_keys_13_1_3, io_keys_13_2_0, io_keys_13_2_1, io_keys_13_2_2, io_keys_13_2_3, io_keys_13_3_0, io_keys_13_3_1, io_keys_13_3_2, io_keys_13_3_3, io_keys_14_0_0, io_keys_14_0_1, io_keys_14_0_2, io_keys_14_0_3, io_keys_14_1_0, io_keys_14_1_1, io_keys_14_1_2, io_keys_14_1_3, io_keys_14_2_0, io_keys_14_2_1, io_keys_14_2_2, io_keys_14_2_3, io_keys_14_3_0, io_keys_14_3_1, io_keys_14_3_2, io_keys_14_3_3, io_aes256, io_shiftCyc, io_shiftRev, io_shift, io_ready, io_dataOut, io_ivOut, io_outputValid);
  (* src = "crypto_accelerator.v:6247" *)
  wire [127:0] _0000_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0001_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0002_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0003_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0004_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0005_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0006_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0007_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0008_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0009_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0010_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0011_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0012_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0013_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0014_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0015_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [7:0] _0016_;
  (* src = "crypto_accelerator.v:6247" *)
  wire [5:0] _0017_;
  (* src = "crypto_accelerator.v:5819" *)
  wire _0018_;
  (* src = "crypto_accelerator.v:5835" *)
  wire _0019_;
  (* src = "crypto_accelerator.v:5851" *)
  wire _0020_;
  (* src = "crypto_accelerator.v:5867" *)
  wire _0021_;
  (* src = "crypto_accelerator.v:5883" *)
  wire _0022_;
  (* src = "crypto_accelerator.v:5899" *)
  wire _0023_;
  (* src = "crypto_accelerator.v:5915" *)
  wire _0024_;
  wire [7:0] _0025_;
  wire [7:0] _0026_;
  wire [7:0] _0027_;
  wire [7:0] _0028_;
  wire [7:0] _0029_;
  wire [7:0] _0030_;
  wire [7:0] _0031_;
  wire [7:0] _0032_;
  wire [7:0] _0033_;
  wire [7:0] _0034_;
  wire [7:0] _0035_;
  wire [7:0] _0036_;
  wire [7:0] _0037_;
  wire [7:0] _0038_;
  wire [7:0] _0039_;
  wire [7:0] _0040_;
  wire [7:0] _0041_;
  wire [7:0] _0042_;
  wire [7:0] _0043_;
  wire [7:0] _0044_;
  wire [7:0] _0045_;
  wire [7:0] _0046_;
  wire [7:0] _0047_;
  wire [7:0] _0048_;
  wire [7:0] _0049_;
  wire [7:0] _0050_;
  wire [7:0] _0051_;
  wire [7:0] _0052_;
  wire [7:0] _0053_;
  wire [7:0] _0054_;
  wire [7:0] _0055_;
  wire [7:0] _0056_;
  wire [7:0] _0057_;
  wire [7:0] _0058_;
  wire [7:0] _0059_;
  wire [7:0] _0060_;
  wire [7:0] _0061_;
  wire [7:0] _0062_;
  wire [7:0] _0063_;
  wire [7:0] _0064_;
  wire [7:0] _0065_;
  wire [7:0] _0066_;
  wire [7:0] _0067_;
  wire [7:0] _0068_;
  wire [7:0] _0069_;
  wire [7:0] _0070_;
  wire [7:0] _0071_;
  wire [7:0] _0072_;
  wire [7:0] _0073_;
  wire [7:0] _0074_;
  wire [7:0] _0075_;
  wire [7:0] _0076_;
  wire [7:0] _0077_;
  wire [7:0] _0078_;
  wire [7:0] _0079_;
  wire [7:0] _0080_;
  wire [7:0] _0081_;
  wire [7:0] _0082_;
  wire [7:0] _0083_;
  wire [7:0] _0084_;
  wire [7:0] _0085_;
  wire [7:0] _0086_;
  wire [7:0] _0087_;
  wire [7:0] _0088_;
  wire [5:0] _0089_;
  wire [5:0] _0090_;
  (* src = "crypto_accelerator.v:3444" *)
  wire [7:0] MixColsModule_io_in_0_0;
  (* src = "crypto_accelerator.v:3445" *)
  wire [7:0] MixColsModule_io_in_0_1;
  (* src = "crypto_accelerator.v:3446" *)
  wire [7:0] MixColsModule_io_in_0_2;
  (* src = "crypto_accelerator.v:3447" *)
  wire [7:0] MixColsModule_io_in_0_3;
  (* src = "crypto_accelerator.v:3448" *)
  wire [7:0] MixColsModule_io_in_1_0;
  (* src = "crypto_accelerator.v:3449" *)
  wire [7:0] MixColsModule_io_in_1_1;
  (* src = "crypto_accelerator.v:3450" *)
  wire [7:0] MixColsModule_io_in_1_2;
  (* src = "crypto_accelerator.v:3451" *)
  wire [7:0] MixColsModule_io_in_1_3;
  (* src = "crypto_accelerator.v:3452" *)
  wire [7:0] MixColsModule_io_in_2_0;
  (* src = "crypto_accelerator.v:3453" *)
  wire [7:0] MixColsModule_io_in_2_1;
  (* src = "crypto_accelerator.v:3454" *)
  wire [7:0] MixColsModule_io_in_2_2;
  (* src = "crypto_accelerator.v:3455" *)
  wire [7:0] MixColsModule_io_in_2_3;
  (* src = "crypto_accelerator.v:3456" *)
  wire [7:0] MixColsModule_io_in_3_0;
  (* src = "crypto_accelerator.v:3457" *)
  wire [7:0] MixColsModule_io_in_3_1;
  (* src = "crypto_accelerator.v:3458" *)
  wire [7:0] MixColsModule_io_in_3_2;
  (* src = "crypto_accelerator.v:3459" *)
  wire [7:0] MixColsModule_io_in_3_3;
  (* src = "crypto_accelerator.v:3460" *)
  wire [7:0] MixColsModule_io_out_0_0;
  (* src = "crypto_accelerator.v:3461" *)
  wire [7:0] MixColsModule_io_out_0_1;
  (* src = "crypto_accelerator.v:3462" *)
  wire [7:0] MixColsModule_io_out_0_2;
  (* src = "crypto_accelerator.v:3463" *)
  wire [7:0] MixColsModule_io_out_0_3;
  (* src = "crypto_accelerator.v:3464" *)
  wire [7:0] MixColsModule_io_out_1_0;
  (* src = "crypto_accelerator.v:3465" *)
  wire [7:0] MixColsModule_io_out_1_1;
  (* src = "crypto_accelerator.v:3466" *)
  wire [7:0] MixColsModule_io_out_1_2;
  (* src = "crypto_accelerator.v:3467" *)
  wire [7:0] MixColsModule_io_out_1_3;
  (* src = "crypto_accelerator.v:3468" *)
  wire [7:0] MixColsModule_io_out_2_0;
  (* src = "crypto_accelerator.v:3469" *)
  wire [7:0] MixColsModule_io_out_2_1;
  (* src = "crypto_accelerator.v:3470" *)
  wire [7:0] MixColsModule_io_out_2_2;
  (* src = "crypto_accelerator.v:3471" *)
  wire [7:0] MixColsModule_io_out_2_3;
  (* src = "crypto_accelerator.v:3472" *)
  wire [7:0] MixColsModule_io_out_3_0;
  (* src = "crypto_accelerator.v:3473" *)
  wire [7:0] MixColsModule_io_out_3_1;
  (* src = "crypto_accelerator.v:3474" *)
  wire [7:0] MixColsModule_io_out_3_2;
  (* src = "crypto_accelerator.v:3475" *)
  wire [7:0] MixColsModule_io_out_3_3;
  (* src = "crypto_accelerator.v:5791" *)
  wire [7:0] _GEN_100;
  (* src = "crypto_accelerator.v:5792" *)
  wire [7:0] _GEN_101;
  (* src = "crypto_accelerator.v:5793" *)
  wire [7:0] _GEN_102;
  (* src = "crypto_accelerator.v:5794" *)
  wire [7:0] _GEN_103;
  (* src = "crypto_accelerator.v:5795" *)
  wire [7:0] _GEN_104;
  (* src = "crypto_accelerator.v:5796" *)
  wire [7:0] _GEN_105;
  (* src = "crypto_accelerator.v:5797" *)
  wire [7:0] _GEN_106;
  (* src = "crypto_accelerator.v:5798" *)
  wire [7:0] _GEN_107;
  (* src = "crypto_accelerator.v:5799" *)
  wire [7:0] _GEN_108;
  (* src = "crypto_accelerator.v:5800" *)
  wire [7:0] _GEN_109;
  (* src = "crypto_accelerator.v:5801" *)
  wire [7:0] _GEN_110;
  (* src = "crypto_accelerator.v:5802" *)
  wire [7:0] _GEN_111;
  (* src = "crypto_accelerator.v:5803" *)
  wire [7:0] _GEN_112;
  (* src = "crypto_accelerator.v:5804" *)
  wire [7:0] _GEN_113;
  (* src = "crypto_accelerator.v:5805" *)
  wire [7:0] _GEN_114;
  (* src = "crypto_accelerator.v:5806" *)
  wire [7:0] _GEN_115;
  (* src = "crypto_accelerator.v:5807" *)
  wire [7:0] _GEN_116;
  (* src = "crypto_accelerator.v:5808" *)
  wire [7:0] _GEN_117;
  (* src = "crypto_accelerator.v:5809" *)
  wire [7:0] _GEN_118;
  (* src = "crypto_accelerator.v:5810" *)
  wire [7:0] _GEN_119;
  (* src = "crypto_accelerator.v:5811" *)
  wire [7:0] _GEN_120;
  (* src = "crypto_accelerator.v:5812" *)
  wire [7:0] _GEN_121;
  (* src = "crypto_accelerator.v:5813" *)
  wire [7:0] _GEN_122;
  (* src = "crypto_accelerator.v:5814" *)
  wire [7:0] _GEN_123;
  (* src = "crypto_accelerator.v:5815" *)
  wire [7:0] _GEN_124;
  (* src = "crypto_accelerator.v:5816" *)
  wire [7:0] _GEN_125;
  (* src = "crypto_accelerator.v:5817" *)
  wire [7:0] _GEN_126;
  (* src = "crypto_accelerator.v:5818" *)
  wire [7:0] _GEN_127;
  (* src = "crypto_accelerator.v:5819" *)
  wire [7:0] _GEN_128;
  (* src = "crypto_accelerator.v:5820" *)
  wire [7:0] _GEN_129;
  (* src = "crypto_accelerator.v:5821" *)
  wire [7:0] _GEN_130;
  (* src = "crypto_accelerator.v:5822" *)
  wire [7:0] _GEN_131;
  (* src = "crypto_accelerator.v:5823" *)
  wire [7:0] _GEN_132;
  (* src = "crypto_accelerator.v:5824" *)
  wire [7:0] _GEN_133;
  (* src = "crypto_accelerator.v:5825" *)
  wire [7:0] _GEN_134;
  (* src = "crypto_accelerator.v:5826" *)
  wire [7:0] _GEN_135;
  (* src = "crypto_accelerator.v:5827" *)
  wire [7:0] _GEN_136;
  (* src = "crypto_accelerator.v:5828" *)
  wire [7:0] _GEN_137;
  (* src = "crypto_accelerator.v:5829" *)
  wire [7:0] _GEN_138;
  (* src = "crypto_accelerator.v:5830" *)
  wire [7:0] _GEN_139;
  (* src = "crypto_accelerator.v:5831" *)
  wire [7:0] _GEN_140;
  (* src = "crypto_accelerator.v:5832" *)
  wire [7:0] _GEN_141;
  (* src = "crypto_accelerator.v:5833" *)
  wire [7:0] _GEN_142;
  (* src = "crypto_accelerator.v:5834" *)
  wire [7:0] _GEN_143;
  (* src = "crypto_accelerator.v:5835" *)
  wire [7:0] _GEN_144;
  (* src = "crypto_accelerator.v:5836" *)
  wire [7:0] _GEN_145;
  (* src = "crypto_accelerator.v:5837" *)
  wire [7:0] _GEN_146;
  (* src = "crypto_accelerator.v:5838" *)
  wire [7:0] _GEN_147;
  (* src = "crypto_accelerator.v:5839" *)
  wire [7:0] _GEN_148;
  (* src = "crypto_accelerator.v:5840" *)
  wire [7:0] _GEN_149;
  (* src = "crypto_accelerator.v:5841" *)
  wire [7:0] _GEN_150;
  (* src = "crypto_accelerator.v:5842" *)
  wire [7:0] _GEN_151;
  (* src = "crypto_accelerator.v:5843" *)
  wire [7:0] _GEN_152;
  (* src = "crypto_accelerator.v:5844" *)
  wire [7:0] _GEN_153;
  (* src = "crypto_accelerator.v:5845" *)
  wire [7:0] _GEN_154;
  (* src = "crypto_accelerator.v:5846" *)
  wire [7:0] _GEN_155;
  (* src = "crypto_accelerator.v:5847" *)
  wire [7:0] _GEN_156;
  (* src = "crypto_accelerator.v:5848" *)
  wire [7:0] _GEN_157;
  (* src = "crypto_accelerator.v:5849" *)
  wire [7:0] _GEN_158;
  (* src = "crypto_accelerator.v:5850" *)
  wire [7:0] _GEN_159;
  (* src = "crypto_accelerator.v:5707" *)
  wire [7:0] _GEN_16;
  (* src = "crypto_accelerator.v:5851" *)
  wire [7:0] _GEN_160;
  (* src = "crypto_accelerator.v:5852" *)
  wire [7:0] _GEN_161;
  (* src = "crypto_accelerator.v:5853" *)
  wire [7:0] _GEN_162;
  (* src = "crypto_accelerator.v:5854" *)
  wire [7:0] _GEN_163;
  (* src = "crypto_accelerator.v:5855" *)
  wire [7:0] _GEN_164;
  (* src = "crypto_accelerator.v:5856" *)
  wire [7:0] _GEN_165;
  (* src = "crypto_accelerator.v:5857" *)
  wire [7:0] _GEN_166;
  (* src = "crypto_accelerator.v:5858" *)
  wire [7:0] _GEN_167;
  (* src = "crypto_accelerator.v:5859" *)
  wire [7:0] _GEN_168;
  (* src = "crypto_accelerator.v:5860" *)
  wire [7:0] _GEN_169;
  (* src = "crypto_accelerator.v:5708" *)
  wire [7:0] _GEN_17;
  (* src = "crypto_accelerator.v:5861" *)
  wire [7:0] _GEN_170;
  (* src = "crypto_accelerator.v:5862" *)
  wire [7:0] _GEN_171;
  (* src = "crypto_accelerator.v:5863" *)
  wire [7:0] _GEN_172;
  (* src = "crypto_accelerator.v:5864" *)
  wire [7:0] _GEN_173;
  (* src = "crypto_accelerator.v:5865" *)
  wire [7:0] _GEN_174;
  (* src = "crypto_accelerator.v:5866" *)
  wire [7:0] _GEN_175;
  (* src = "crypto_accelerator.v:5867" *)
  wire [7:0] _GEN_176;
  (* src = "crypto_accelerator.v:5868" *)
  wire [7:0] _GEN_177;
  (* src = "crypto_accelerator.v:5869" *)
  wire [7:0] _GEN_178;
  (* src = "crypto_accelerator.v:5870" *)
  wire [7:0] _GEN_179;
  (* src = "crypto_accelerator.v:5709" *)
  wire [7:0] _GEN_18;
  (* src = "crypto_accelerator.v:5871" *)
  wire [7:0] _GEN_180;
  (* src = "crypto_accelerator.v:5872" *)
  wire [7:0] _GEN_181;
  (* src = "crypto_accelerator.v:5873" *)
  wire [7:0] _GEN_182;
  (* src = "crypto_accelerator.v:5874" *)
  wire [7:0] _GEN_183;
  (* src = "crypto_accelerator.v:5875" *)
  wire [7:0] _GEN_184;
  (* src = "crypto_accelerator.v:5876" *)
  wire [7:0] _GEN_185;
  (* src = "crypto_accelerator.v:5877" *)
  wire [7:0] _GEN_186;
  (* src = "crypto_accelerator.v:5878" *)
  wire [7:0] _GEN_187;
  (* src = "crypto_accelerator.v:5879" *)
  wire [7:0] _GEN_188;
  (* src = "crypto_accelerator.v:5880" *)
  wire [7:0] _GEN_189;
  (* src = "crypto_accelerator.v:5710" *)
  wire [7:0] _GEN_19;
  (* src = "crypto_accelerator.v:5881" *)
  wire [7:0] _GEN_190;
  (* src = "crypto_accelerator.v:5882" *)
  wire [7:0] _GEN_191;
  (* src = "crypto_accelerator.v:5883" *)
  wire [7:0] _GEN_192;
  (* src = "crypto_accelerator.v:5884" *)
  wire [7:0] _GEN_193;
  (* src = "crypto_accelerator.v:5885" *)
  wire [7:0] _GEN_194;
  (* src = "crypto_accelerator.v:5886" *)
  wire [7:0] _GEN_195;
  (* src = "crypto_accelerator.v:5887" *)
  wire [7:0] _GEN_196;
  (* src = "crypto_accelerator.v:5888" *)
  wire [7:0] _GEN_197;
  (* src = "crypto_accelerator.v:5889" *)
  wire [7:0] _GEN_198;
  (* src = "crypto_accelerator.v:5890" *)
  wire [7:0] _GEN_199;
  (* src = "crypto_accelerator.v:5711" *)
  wire [7:0] _GEN_20;
  (* src = "crypto_accelerator.v:5891" *)
  wire [7:0] _GEN_200;
  (* src = "crypto_accelerator.v:5892" *)
  wire [7:0] _GEN_201;
  (* src = "crypto_accelerator.v:5893" *)
  wire [7:0] _GEN_202;
  (* src = "crypto_accelerator.v:5894" *)
  wire [7:0] _GEN_203;
  (* src = "crypto_accelerator.v:5895" *)
  wire [7:0] _GEN_204;
  (* src = "crypto_accelerator.v:5896" *)
  wire [7:0] _GEN_205;
  (* src = "crypto_accelerator.v:5897" *)
  wire [7:0] _GEN_206;
  (* src = "crypto_accelerator.v:5898" *)
  wire [7:0] _GEN_207;
  (* src = "crypto_accelerator.v:5899" *)
  wire [7:0] _GEN_208;
  (* src = "crypto_accelerator.v:5900" *)
  wire [7:0] _GEN_209;
  (* src = "crypto_accelerator.v:5712" *)
  wire [7:0] _GEN_21;
  (* src = "crypto_accelerator.v:5901" *)
  wire [7:0] _GEN_210;
  (* src = "crypto_accelerator.v:5902" *)
  wire [7:0] _GEN_211;
  (* src = "crypto_accelerator.v:5903" *)
  wire [7:0] _GEN_212;
  (* src = "crypto_accelerator.v:5904" *)
  wire [7:0] _GEN_213;
  (* src = "crypto_accelerator.v:5905" *)
  wire [7:0] _GEN_214;
  (* src = "crypto_accelerator.v:5906" *)
  wire [7:0] _GEN_215;
  (* src = "crypto_accelerator.v:5907" *)
  wire [7:0] _GEN_216;
  (* src = "crypto_accelerator.v:5908" *)
  wire [7:0] _GEN_217;
  (* src = "crypto_accelerator.v:5909" *)
  wire [7:0] _GEN_218;
  (* src = "crypto_accelerator.v:5910" *)
  wire [7:0] _GEN_219;
  (* src = "crypto_accelerator.v:5713" *)
  wire [7:0] _GEN_22;
  (* src = "crypto_accelerator.v:5911" *)
  wire [7:0] _GEN_220;
  (* src = "crypto_accelerator.v:5912" *)
  wire [7:0] _GEN_221;
  (* src = "crypto_accelerator.v:5913" *)
  wire [7:0] _GEN_222;
  (* src = "crypto_accelerator.v:5914" *)
  wire [7:0] _GEN_223;
  (* src = "crypto_accelerator.v:5915" *)
  wire [7:0] _GEN_224;
  (* src = "crypto_accelerator.v:5916" *)
  wire [7:0] _GEN_225;
  (* src = "crypto_accelerator.v:5917" *)
  wire [7:0] _GEN_226;
  (* src = "crypto_accelerator.v:5918" *)
  wire [7:0] _GEN_227;
  (* src = "crypto_accelerator.v:5919" *)
  wire [7:0] _GEN_228;
  (* src = "crypto_accelerator.v:5920" *)
  wire [7:0] _GEN_229;
  (* src = "crypto_accelerator.v:5714" *)
  wire [7:0] _GEN_23;
  (* src = "crypto_accelerator.v:5921" *)
  wire [7:0] _GEN_230;
  (* src = "crypto_accelerator.v:5922" *)
  wire [7:0] _GEN_231;
  (* src = "crypto_accelerator.v:5923" *)
  wire [7:0] _GEN_232;
  (* src = "crypto_accelerator.v:5924" *)
  wire [7:0] _GEN_233;
  (* src = "crypto_accelerator.v:5925" *)
  wire [7:0] _GEN_234;
  (* src = "crypto_accelerator.v:5926" *)
  wire [7:0] _GEN_235;
  (* src = "crypto_accelerator.v:5927" *)
  wire [7:0] _GEN_236;
  (* src = "crypto_accelerator.v:5928" *)
  wire [7:0] _GEN_237;
  (* src = "crypto_accelerator.v:5929" *)
  wire [7:0] _GEN_238;
  (* src = "crypto_accelerator.v:5930" *)
  wire [7:0] _GEN_239;
  (* src = "crypto_accelerator.v:5715" *)
  wire [7:0] _GEN_24;
  (* src = "crypto_accelerator.v:5716" *)
  wire [7:0] _GEN_25;
  (* src = "crypto_accelerator.v:5717" *)
  wire [7:0] _GEN_26;
  (* src = "crypto_accelerator.v:5718" *)
  wire [7:0] _GEN_27;
  (* src = "crypto_accelerator.v:6109" *)
  wire _GEN_275;
  (* src = "crypto_accelerator.v:5719" *)
  wire [7:0] _GEN_28;
  (* src = "crypto_accelerator.v:5720" *)
  wire [7:0] _GEN_29;
  (* src = "crypto_accelerator.v:6110" *)
  wire _GEN_292;
  (* src = "crypto_accelerator.v:5721" *)
  wire [7:0] _GEN_30;
  (* src = "crypto_accelerator.v:5722" *)
  wire [7:0] _GEN_31;
  (* src = "crypto_accelerator.v:5973" *)
  wire [9:0] _GEN_311;
  (* src = "crypto_accelerator.v:5975" *)
  wire [9:0] _GEN_312;
  (* src = "crypto_accelerator.v:5977" *)
  wire [9:0] _GEN_313;
  (* src = "crypto_accelerator.v:5979" *)
  wire [9:0] _GEN_314;
  (* src = "crypto_accelerator.v:6007" *)
  wire [9:0] _GEN_315;
  (* src = "crypto_accelerator.v:6009" *)
  wire [9:0] _GEN_316;
  (* src = "crypto_accelerator.v:6011" *)
  wire [9:0] _GEN_317;
  (* src = "crypto_accelerator.v:6013" *)
  wire [9:0] _GEN_318;
  (* src = "crypto_accelerator.v:6041" *)
  wire [9:0] _GEN_319;
  (* src = "crypto_accelerator.v:5723" *)
  wire [7:0] _GEN_32;
  (* src = "crypto_accelerator.v:6043" *)
  wire [9:0] _GEN_320;
  (* src = "crypto_accelerator.v:6045" *)
  wire [9:0] _GEN_321;
  (* src = "crypto_accelerator.v:6047" *)
  wire [9:0] _GEN_322;
  (* src = "crypto_accelerator.v:6075" *)
  wire [9:0] _GEN_323;
  (* src = "crypto_accelerator.v:6077" *)
  wire [9:0] _GEN_324;
  (* src = "crypto_accelerator.v:6079" *)
  wire [9:0] _GEN_325;
  (* src = "crypto_accelerator.v:6081" *)
  wire [9:0] _GEN_326;
  wire [3:0] _GEN_327;
  (* src = "crypto_accelerator.v:5724" *)
  wire [7:0] _GEN_33;
  (* src = "crypto_accelerator.v:5725" *)
  wire [7:0] _GEN_34;
  (* src = "crypto_accelerator.v:5726" *)
  wire [7:0] _GEN_35;
  (* src = "crypto_accelerator.v:5727" *)
  wire [7:0] _GEN_36;
  (* src = "crypto_accelerator.v:5728" *)
  wire [7:0] _GEN_37;
  (* src = "crypto_accelerator.v:5729" *)
  wire [7:0] _GEN_38;
  (* src = "crypto_accelerator.v:5730" *)
  wire [7:0] _GEN_39;
  (* src = "crypto_accelerator.v:5731" *)
  wire [7:0] _GEN_40;
  (* src = "crypto_accelerator.v:5732" *)
  wire [7:0] _GEN_41;
  (* src = "crypto_accelerator.v:5733" *)
  wire [7:0] _GEN_42;
  (* src = "crypto_accelerator.v:5734" *)
  wire [7:0] _GEN_43;
  (* src = "crypto_accelerator.v:5735" *)
  wire [7:0] _GEN_44;
  (* src = "crypto_accelerator.v:5736" *)
  wire [7:0] _GEN_45;
  (* src = "crypto_accelerator.v:5737" *)
  wire [7:0] _GEN_46;
  (* src = "crypto_accelerator.v:5738" *)
  wire [7:0] _GEN_47;
  (* src = "crypto_accelerator.v:5739" *)
  wire [7:0] _GEN_48;
  (* src = "crypto_accelerator.v:5740" *)
  wire [7:0] _GEN_49;
  (* src = "crypto_accelerator.v:5741" *)
  wire [7:0] _GEN_50;
  (* src = "crypto_accelerator.v:5742" *)
  wire [7:0] _GEN_51;
  (* src = "crypto_accelerator.v:5743" *)
  wire [7:0] _GEN_52;
  (* src = "crypto_accelerator.v:5744" *)
  wire [7:0] _GEN_53;
  (* src = "crypto_accelerator.v:5745" *)
  wire [7:0] _GEN_54;
  (* src = "crypto_accelerator.v:5746" *)
  wire [7:0] _GEN_55;
  (* src = "crypto_accelerator.v:5747" *)
  wire [7:0] _GEN_56;
  (* src = "crypto_accelerator.v:5748" *)
  wire [7:0] _GEN_57;
  (* src = "crypto_accelerator.v:5749" *)
  wire [7:0] _GEN_58;
  (* src = "crypto_accelerator.v:5750" *)
  wire [7:0] _GEN_59;
  (* src = "crypto_accelerator.v:5751" *)
  wire [7:0] _GEN_60;
  (* src = "crypto_accelerator.v:5752" *)
  wire [7:0] _GEN_61;
  (* src = "crypto_accelerator.v:5753" *)
  wire [7:0] _GEN_62;
  (* src = "crypto_accelerator.v:5754" *)
  wire [7:0] _GEN_63;
  (* src = "crypto_accelerator.v:5755" *)
  wire [7:0] _GEN_64;
  (* src = "crypto_accelerator.v:5756" *)
  wire [7:0] _GEN_65;
  (* src = "crypto_accelerator.v:5757" *)
  wire [7:0] _GEN_66;
  (* src = "crypto_accelerator.v:5758" *)
  wire [7:0] _GEN_67;
  (* src = "crypto_accelerator.v:5759" *)
  wire [7:0] _GEN_68;
  (* src = "crypto_accelerator.v:5760" *)
  wire [7:0] _GEN_69;
  (* src = "crypto_accelerator.v:5761" *)
  wire [7:0] _GEN_70;
  (* src = "crypto_accelerator.v:5762" *)
  wire [7:0] _GEN_71;
  (* src = "crypto_accelerator.v:5763" *)
  wire [7:0] _GEN_72;
  (* src = "crypto_accelerator.v:5764" *)
  wire [7:0] _GEN_73;
  (* src = "crypto_accelerator.v:5765" *)
  wire [7:0] _GEN_74;
  (* src = "crypto_accelerator.v:5766" *)
  wire [7:0] _GEN_75;
  (* src = "crypto_accelerator.v:5767" *)
  wire [7:0] _GEN_76;
  (* src = "crypto_accelerator.v:5768" *)
  wire [7:0] _GEN_77;
  (* src = "crypto_accelerator.v:5769" *)
  wire [7:0] _GEN_78;
  (* src = "crypto_accelerator.v:5770" *)
  wire [7:0] _GEN_79;
  (* src = "crypto_accelerator.v:5771" *)
  wire [7:0] _GEN_80;
  (* src = "crypto_accelerator.v:5772" *)
  wire [7:0] _GEN_81;
  (* src = "crypto_accelerator.v:5773" *)
  wire [7:0] _GEN_82;
  (* src = "crypto_accelerator.v:5774" *)
  wire [7:0] _GEN_83;
  (* src = "crypto_accelerator.v:5775" *)
  wire [7:0] _GEN_84;
  (* src = "crypto_accelerator.v:5776" *)
  wire [7:0] _GEN_85;
  (* src = "crypto_accelerator.v:5777" *)
  wire [7:0] _GEN_86;
  (* src = "crypto_accelerator.v:5778" *)
  wire [7:0] _GEN_87;
  (* src = "crypto_accelerator.v:5779" *)
  wire [7:0] _GEN_88;
  (* src = "crypto_accelerator.v:5780" *)
  wire [7:0] _GEN_89;
  (* src = "crypto_accelerator.v:5781" *)
  wire [7:0] _GEN_90;
  (* src = "crypto_accelerator.v:5782" *)
  wire [7:0] _GEN_91;
  (* src = "crypto_accelerator.v:5783" *)
  wire [7:0] _GEN_92;
  (* src = "crypto_accelerator.v:5784" *)
  wire [7:0] _GEN_93;
  (* src = "crypto_accelerator.v:5785" *)
  wire [7:0] _GEN_94;
  (* src = "crypto_accelerator.v:5786" *)
  wire [7:0] _GEN_95;
  (* src = "crypto_accelerator.v:5787" *)
  wire [7:0] _GEN_96;
  (* src = "crypto_accelerator.v:5788" *)
  wire [7:0] _GEN_97;
  (* src = "crypto_accelerator.v:5789" *)
  wire [7:0] _GEN_98;
  (* src = "crypto_accelerator.v:5790" *)
  wire [7:0] _GEN_99;
  (* src = "crypto_accelerator.v:3477" *)
  wire _T;
  (* src = "crypto_accelerator.v:3478" *)
  wire _T_1;
  (* src = "crypto_accelerator.v:3496" *)
  wire [63:0] _T_10;
  (* src = "crypto_accelerator.v:3978" *)
  wire _T_1000;
  (* src = "crypto_accelerator.v:3979" *)
  wire _T_1002;
  (* src = "crypto_accelerator.v:3980" *)
  wire _T_1004;
  (* src = "crypto_accelerator.v:3981" *)
  wire _T_1006;
  (* src = "crypto_accelerator.v:3982" *)
  wire _T_1008;
  (* src = "crypto_accelerator.v:3533" *)
  wire _T_101;
  (* src = "crypto_accelerator.v:3983" *)
  wire _T_1010;
  (* src = "crypto_accelerator.v:3984" *)
  wire _T_1012;
  (* src = "crypto_accelerator.v:3985" *)
  wire _T_1014;
  (* src = "crypto_accelerator.v:3986" *)
  wire _T_1016;
  (* src = "crypto_accelerator.v:3987" *)
  wire _T_1018;
  (* src = "crypto_accelerator.v:3988" *)
  wire _T_1020;
  (* src = "crypto_accelerator.v:3989" *)
  wire _T_1022;
  (* src = "crypto_accelerator.v:3990" *)
  wire _T_1024;
  (* src = "crypto_accelerator.v:3991" *)
  wire _T_1026;
  (* src = "crypto_accelerator.v:3992" *)
  wire _T_1028;
  (* src = "crypto_accelerator.v:3534" *)
  wire _T_103;
  (* src = "crypto_accelerator.v:3993" *)
  wire _T_1030;
  (* src = "crypto_accelerator.v:3994" *)
  wire _T_1032;
  (* src = "crypto_accelerator.v:3995" *)
  wire _T_1034;
  (* src = "crypto_accelerator.v:3996" *)
  wire _T_1036;
  (* src = "crypto_accelerator.v:3997" *)
  wire _T_1038;
  (* src = "crypto_accelerator.v:3998" *)
  wire _T_1040;
  (* src = "crypto_accelerator.v:3999" *)
  wire _T_1042;
  (* src = "crypto_accelerator.v:4000" *)
  wire _T_1044;
  (* src = "crypto_accelerator.v:4001" *)
  wire _T_1046;
  (* src = "crypto_accelerator.v:4002" *)
  wire _T_1048;
  (* src = "crypto_accelerator.v:3535" *)
  wire _T_105;
  (* src = "crypto_accelerator.v:4003" *)
  wire _T_1050;
  (* src = "crypto_accelerator.v:4004" *)
  wire _T_1052;
  (* src = "crypto_accelerator.v:4005" *)
  wire _T_1054;
  (* src = "crypto_accelerator.v:4006" *)
  wire _T_1056;
  (* src = "crypto_accelerator.v:4007" *)
  wire _T_1058;
  (* src = "crypto_accelerator.v:4008" *)
  wire _T_1060;
  (* src = "crypto_accelerator.v:4009" *)
  wire _T_1062;
  (* src = "crypto_accelerator.v:4010" *)
  wire _T_1064;
  (* src = "crypto_accelerator.v:4011" *)
  wire _T_1066;
  (* src = "crypto_accelerator.v:4012" *)
  wire _T_1068;
  (* src = "crypto_accelerator.v:3536" *)
  wire _T_107;
  (* src = "crypto_accelerator.v:4013" *)
  wire _T_1070;
  (* src = "crypto_accelerator.v:4014" *)
  wire _T_1072;
  (* src = "crypto_accelerator.v:4015" *)
  wire _T_1074;
  (* src = "crypto_accelerator.v:4016" *)
  wire _T_1076;
  (* src = "crypto_accelerator.v:4017" *)
  wire _T_1078;
  (* src = "crypto_accelerator.v:4018" *)
  wire _T_1080;
  (* src = "crypto_accelerator.v:4019" *)
  wire _T_1082;
  (* src = "crypto_accelerator.v:4020" *)
  wire _T_1084;
  (* src = "crypto_accelerator.v:4021" *)
  wire _T_1086;
  (* src = "crypto_accelerator.v:4022" *)
  wire _T_1088;
  (* src = "crypto_accelerator.v:3537" *)
  wire _T_109;
  (* src = "crypto_accelerator.v:4023" *)
  wire _T_1090;
  (* src = "crypto_accelerator.v:4024" *)
  wire _T_1092;
  (* src = "crypto_accelerator.v:4025" *)
  wire _T_1094;
  (* src = "crypto_accelerator.v:4026" *)
  wire _T_1096;
  (* src = "crypto_accelerator.v:4027" *)
  wire _T_1098;
  (* src = "crypto_accelerator.v:4028" *)
  wire _T_1100;
  (* src = "crypto_accelerator.v:4029" *)
  wire _T_1102;
  (* src = "crypto_accelerator.v:4030" *)
  wire _T_1104;
  (* src = "crypto_accelerator.v:4031" *)
  wire _T_1106;
  (* src = "crypto_accelerator.v:4032" *)
  wire _T_1108;
  (* src = "crypto_accelerator.v:3538" *)
  wire _T_111;
  (* src = "crypto_accelerator.v:4033" *)
  wire _T_1110;
  (* src = "crypto_accelerator.v:4034" *)
  wire _T_1112;
  (* src = "crypto_accelerator.v:4035" *)
  wire _T_1114;
  (* src = "crypto_accelerator.v:4036" *)
  wire _T_1116;
  (* src = "crypto_accelerator.v:4037" *)
  wire _T_1118;
  (* src = "crypto_accelerator.v:4038" *)
  wire _T_1120;
  (* src = "crypto_accelerator.v:4039" *)
  wire _T_1122;
  (* src = "crypto_accelerator.v:4040" *)
  wire _T_1124;
  (* src = "crypto_accelerator.v:4041" *)
  wire _T_1125;
  (* src = "crypto_accelerator.v:4042" *)
  wire _T_1126;
  (* src = "crypto_accelerator.v:4043" *)
  wire _T_1127;
  (* src = "crypto_accelerator.v:4044" *)
  wire _T_1128;
  (* src = "crypto_accelerator.v:4045" *)
  wire _T_1129;
  (* src = "crypto_accelerator.v:3539" *)
  wire _T_113;
  (* src = "crypto_accelerator.v:4046" *)
  wire _T_1130;
  (* src = "crypto_accelerator.v:4047" *)
  wire _T_1131;
  (* src = "crypto_accelerator.v:4048" *)
  wire _T_1132;
  (* src = "crypto_accelerator.v:3540" *)
  wire _T_115;
  (* src = "crypto_accelerator.v:4050" *)
  wire _T_1158;
  (* src = "crypto_accelerator.v:4051" *)
  wire _T_1160;
  (* src = "crypto_accelerator.v:4052" *)
  wire _T_1161;
  (* src = "crypto_accelerator.v:4053" *)
  wire _T_1163;
  (* src = "crypto_accelerator.v:4054" *)
  wire _T_1164;
  (* src = "crypto_accelerator.v:4055" *)
  wire _T_1166;
  (* src = "crypto_accelerator.v:4056" *)
  wire _T_1168;
  (* src = "crypto_accelerator.v:4057" *)
  wire _T_1169;
  (* src = "crypto_accelerator.v:3541" *)
  wire _T_117;
  (* src = "crypto_accelerator.v:4058" *)
  wire _T_1171;
  (* src = "crypto_accelerator.v:4059" *)
  wire _T_1173;
  (* src = "crypto_accelerator.v:4060" *)
  wire _T_1174;
  (* src = "crypto_accelerator.v:4061" *)
  wire _T_1176;
  (* src = "crypto_accelerator.v:4062" *)
  wire _T_1178;
  (* src = "crypto_accelerator.v:4063" *)
  wire _T_1179;
  (* src = "crypto_accelerator.v:4064" *)
  wire _T_1181;
  (* src = "crypto_accelerator.v:4065" *)
  wire _T_1183;
  (* src = "crypto_accelerator.v:4066" *)
  wire _T_1185;
  (* src = "crypto_accelerator.v:4067" *)
  wire _T_1187;
  (* src = "crypto_accelerator.v:4068" *)
  wire _T_1188;
  (* src = "crypto_accelerator.v:3542" *)
  wire _T_119;
  (* src = "crypto_accelerator.v:4069" *)
  wire _T_1190;
  (* src = "crypto_accelerator.v:4070" *)
  wire _T_1192;
  (* src = "crypto_accelerator.v:4071" *)
  wire _T_1193;
  (* src = "crypto_accelerator.v:4072" *)
  wire _T_1195;
  (* src = "crypto_accelerator.v:4073" *)
  wire _T_1197;
  (* src = "crypto_accelerator.v:4074" *)
  wire _T_1199;
  (* src = "crypto_accelerator.v:4075" *)
  wire _T_1200;
  (* src = "crypto_accelerator.v:4076" *)
  wire _T_1202;
  (* src = "crypto_accelerator.v:4077" *)
  wire _T_1203;
  (* src = "crypto_accelerator.v:4078" *)
  wire _T_1205;
  (* src = "crypto_accelerator.v:4079" *)
  wire _T_1206;
  (* src = "crypto_accelerator.v:4080" *)
  wire _T_1208;
  (* src = "crypto_accelerator.v:3543" *)
  wire _T_121;
  (* src = "crypto_accelerator.v:4081" *)
  wire _T_1210;
  (* src = "crypto_accelerator.v:4082" *)
  wire _T_1212;
  (* src = "crypto_accelerator.v:4083" *)
  wire _T_1214;
  (* src = "crypto_accelerator.v:4084" *)
  wire _T_1216;
  (* src = "crypto_accelerator.v:4085" *)
  wire _T_1218;
  (* src = "crypto_accelerator.v:4086" *)
  wire _T_1220;
  (* src = "crypto_accelerator.v:4087" *)
  wire _T_1222;
  (* src = "crypto_accelerator.v:4088" *)
  wire _T_1224;
  (* src = "crypto_accelerator.v:4089" *)
  wire _T_1226;
  (* src = "crypto_accelerator.v:4090" *)
  wire _T_1228;
  (* src = "crypto_accelerator.v:3544" *)
  wire _T_123;
  (* src = "crypto_accelerator.v:4091" *)
  wire _T_1230;
  (* src = "crypto_accelerator.v:4092" *)
  wire _T_1232;
  (* src = "crypto_accelerator.v:4093" *)
  wire _T_1234;
  (* src = "crypto_accelerator.v:4094" *)
  wire _T_1236;
  (* src = "crypto_accelerator.v:4095" *)
  wire _T_1238;
  (* src = "crypto_accelerator.v:4096" *)
  wire _T_1240;
  (* src = "crypto_accelerator.v:4097" *)
  wire _T_1242;
  (* src = "crypto_accelerator.v:4098" *)
  wire _T_1244;
  (* src = "crypto_accelerator.v:4099" *)
  wire _T_1246;
  (* src = "crypto_accelerator.v:4100" *)
  wire _T_1248;
  (* src = "crypto_accelerator.v:3545" *)
  wire _T_125;
  (* src = "crypto_accelerator.v:4101" *)
  wire _T_1250;
  (* src = "crypto_accelerator.v:4102" *)
  wire _T_1252;
  (* src = "crypto_accelerator.v:4103" *)
  wire _T_1254;
  (* src = "crypto_accelerator.v:4104" *)
  wire _T_1256;
  (* src = "crypto_accelerator.v:4105" *)
  wire _T_1258;
  (* src = "crypto_accelerator.v:4106" *)
  wire _T_1260;
  (* src = "crypto_accelerator.v:4107" *)
  wire _T_1262;
  (* src = "crypto_accelerator.v:4108" *)
  wire _T_1264;
  (* src = "crypto_accelerator.v:4109" *)
  wire _T_1266;
  (* src = "crypto_accelerator.v:4110" *)
  wire _T_1268;
  (* src = "crypto_accelerator.v:3546" *)
  wire _T_127;
  (* src = "crypto_accelerator.v:4111" *)
  wire _T_1270;
  (* src = "crypto_accelerator.v:4112" *)
  wire _T_1272;
  (* src = "crypto_accelerator.v:4113" *)
  wire _T_1274;
  (* src = "crypto_accelerator.v:4114" *)
  wire _T_1276;
  (* src = "crypto_accelerator.v:4115" *)
  wire _T_1278;
  (* src = "crypto_accelerator.v:4116" *)
  wire _T_1280;
  (* src = "crypto_accelerator.v:4117" *)
  wire _T_1282;
  (* src = "crypto_accelerator.v:4118" *)
  wire _T_1284;
  (* src = "crypto_accelerator.v:4119" *)
  wire _T_1286;
  (* src = "crypto_accelerator.v:4120" *)
  wire _T_1288;
  (* src = "crypto_accelerator.v:3547" *)
  wire _T_129;
  (* src = "crypto_accelerator.v:4121" *)
  wire _T_1290;
  (* src = "crypto_accelerator.v:4122" *)
  wire _T_1292;
  (* src = "crypto_accelerator.v:4123" *)
  wire _T_1294;
  (* src = "crypto_accelerator.v:4124" *)
  wire _T_1296;
  (* src = "crypto_accelerator.v:4125" *)
  wire _T_1298;
  (* src = "crypto_accelerator.v:4126" *)
  wire _T_1300;
  (* src = "crypto_accelerator.v:4127" *)
  wire _T_1302;
  (* src = "crypto_accelerator.v:4128" *)
  wire _T_1304;
  (* src = "crypto_accelerator.v:4129" *)
  wire _T_1306;
  (* src = "crypto_accelerator.v:4130" *)
  wire _T_1308;
  (* src = "crypto_accelerator.v:3548" *)
  wire _T_131;
  (* src = "crypto_accelerator.v:4131" *)
  wire _T_1310;
  (* src = "crypto_accelerator.v:4132" *)
  wire _T_1312;
  (* src = "crypto_accelerator.v:4133" *)
  wire _T_1314;
  (* src = "crypto_accelerator.v:4134" *)
  wire _T_1316;
  (* src = "crypto_accelerator.v:4135" *)
  wire _T_1318;
  (* src = "crypto_accelerator.v:4136" *)
  wire _T_1320;
  (* src = "crypto_accelerator.v:4137" *)
  wire _T_1322;
  (* src = "crypto_accelerator.v:4138" *)
  wire _T_1324;
  (* src = "crypto_accelerator.v:4139" *)
  wire _T_1326;
  (* src = "crypto_accelerator.v:4140" *)
  wire _T_1328;
  (* src = "crypto_accelerator.v:3549" *)
  wire _T_133;
  (* src = "crypto_accelerator.v:4141" *)
  wire _T_1330;
  (* src = "crypto_accelerator.v:4142" *)
  wire _T_1332;
  (* src = "crypto_accelerator.v:4143" *)
  wire _T_1334;
  (* src = "crypto_accelerator.v:4144" *)
  wire _T_1336;
  (* src = "crypto_accelerator.v:4145" *)
  wire _T_1338;
  (* src = "crypto_accelerator.v:4146" *)
  wire _T_1340;
  (* src = "crypto_accelerator.v:4147" *)
  wire _T_1342;
  (* src = "crypto_accelerator.v:4148" *)
  wire _T_1344;
  (* src = "crypto_accelerator.v:4149" *)
  wire _T_1346;
  (* src = "crypto_accelerator.v:4150" *)
  wire _T_1348;
  (* src = "crypto_accelerator.v:3550" *)
  wire _T_135;
  (* src = "crypto_accelerator.v:4151" *)
  wire _T_1350;
  (* src = "crypto_accelerator.v:4152" *)
  wire _T_1352;
  (* src = "crypto_accelerator.v:4153" *)
  wire _T_1354;
  (* src = "crypto_accelerator.v:4154" *)
  wire _T_1356;
  (* src = "crypto_accelerator.v:4155" *)
  wire _T_1358;
  (* src = "crypto_accelerator.v:4156" *)
  wire _T_1360;
  (* src = "crypto_accelerator.v:4157" *)
  wire _T_1362;
  (* src = "crypto_accelerator.v:4158" *)
  wire _T_1364;
  (* src = "crypto_accelerator.v:4159" *)
  wire _T_1366;
  (* src = "crypto_accelerator.v:4160" *)
  wire _T_1368;
  (* src = "crypto_accelerator.v:3551" *)
  wire _T_137;
  (* src = "crypto_accelerator.v:4161" *)
  wire _T_1370;
  (* src = "crypto_accelerator.v:4162" *)
  wire _T_1372;
  (* src = "crypto_accelerator.v:4163" *)
  wire _T_1374;
  (* src = "crypto_accelerator.v:4164" *)
  wire _T_1376;
  (* src = "crypto_accelerator.v:4165" *)
  wire _T_1378;
  (* src = "crypto_accelerator.v:4166" *)
  wire _T_1380;
  (* src = "crypto_accelerator.v:4167" *)
  wire _T_1382;
  (* src = "crypto_accelerator.v:4168" *)
  wire _T_1384;
  (* src = "crypto_accelerator.v:4169" *)
  wire _T_1386;
  (* src = "crypto_accelerator.v:4170" *)
  wire _T_1388;
  (* src = "crypto_accelerator.v:3552" *)
  wire _T_139;
  (* src = "crypto_accelerator.v:4171" *)
  wire _T_1390;
  (* src = "crypto_accelerator.v:4172" *)
  wire _T_1392;
  (* src = "crypto_accelerator.v:4173" *)
  wire _T_1394;
  (* src = "crypto_accelerator.v:4174" *)
  wire _T_1396;
  (* src = "crypto_accelerator.v:4175" *)
  wire _T_1398;
  (* src = "crypto_accelerator.v:4176" *)
  wire _T_1400;
  (* src = "crypto_accelerator.v:4177" *)
  wire _T_1402;
  (* src = "crypto_accelerator.v:4178" *)
  wire _T_1404;
  (* src = "crypto_accelerator.v:4179" *)
  wire _T_1405;
  (* src = "crypto_accelerator.v:4180" *)
  wire _T_1406;
  (* src = "crypto_accelerator.v:4181" *)
  wire _T_1407;
  (* src = "crypto_accelerator.v:4182" *)
  wire _T_1408;
  (* src = "crypto_accelerator.v:4183" *)
  wire _T_1409;
  (* src = "crypto_accelerator.v:3553" *)
  wire _T_141;
  (* src = "crypto_accelerator.v:4184" *)
  wire _T_1410;
  (* src = "crypto_accelerator.v:4185" *)
  wire _T_1411;
  (* src = "crypto_accelerator.v:4186" *)
  wire _T_1412;
  (* src = "crypto_accelerator.v:3554" *)
  wire _T_143;
  (* src = "crypto_accelerator.v:4188" *)
  wire _T_1437;
  (* src = "crypto_accelerator.v:4189" *)
  wire _T_1439;
  (* src = "crypto_accelerator.v:4190" *)
  wire _T_1440;
  (* src = "crypto_accelerator.v:4191" *)
  wire _T_1442;
  (* src = "crypto_accelerator.v:4192" *)
  wire _T_1443;
  (* src = "crypto_accelerator.v:4193" *)
  wire _T_1445;
  (* src = "crypto_accelerator.v:4194" *)
  wire _T_1447;
  (* src = "crypto_accelerator.v:4195" *)
  wire _T_1448;
  (* src = "crypto_accelerator.v:3555" *)
  wire _T_145;
  (* src = "crypto_accelerator.v:4196" *)
  wire _T_1450;
  (* src = "crypto_accelerator.v:4197" *)
  wire _T_1452;
  (* src = "crypto_accelerator.v:4198" *)
  wire _T_1453;
  (* src = "crypto_accelerator.v:4199" *)
  wire _T_1455;
  (* src = "crypto_accelerator.v:4200" *)
  wire _T_1457;
  (* src = "crypto_accelerator.v:4201" *)
  wire _T_1458;
  (* src = "crypto_accelerator.v:4202" *)
  wire _T_1460;
  (* src = "crypto_accelerator.v:4203" *)
  wire _T_1462;
  (* src = "crypto_accelerator.v:4204" *)
  wire _T_1464;
  (* src = "crypto_accelerator.v:4205" *)
  wire _T_1466;
  (* src = "crypto_accelerator.v:4206" *)
  wire _T_1467;
  (* src = "crypto_accelerator.v:4207" *)
  wire _T_1469;
  (* src = "crypto_accelerator.v:3556" *)
  wire _T_147;
  (* src = "crypto_accelerator.v:4208" *)
  wire _T_1471;
  (* src = "crypto_accelerator.v:4209" *)
  wire _T_1472;
  (* src = "crypto_accelerator.v:4210" *)
  wire _T_1474;
  (* src = "crypto_accelerator.v:4211" *)
  wire _T_1476;
  (* src = "crypto_accelerator.v:4212" *)
  wire _T_1478;
  (* src = "crypto_accelerator.v:4213" *)
  wire _T_1479;
  (* src = "crypto_accelerator.v:4214" *)
  wire _T_1481;
  (* src = "crypto_accelerator.v:4215" *)
  wire _T_1482;
  (* src = "crypto_accelerator.v:4216" *)
  wire _T_1484;
  (* src = "crypto_accelerator.v:4217" *)
  wire _T_1485;
  (* src = "crypto_accelerator.v:4218" *)
  wire _T_1487;
  (* src = "crypto_accelerator.v:4219" *)
  wire _T_1489;
  (* src = "crypto_accelerator.v:3557" *)
  wire _T_149;
  (* src = "crypto_accelerator.v:4220" *)
  wire _T_1491;
  (* src = "crypto_accelerator.v:4221" *)
  wire _T_1493;
  (* src = "crypto_accelerator.v:4222" *)
  wire _T_1495;
  (* src = "crypto_accelerator.v:4223" *)
  wire _T_1497;
  (* src = "crypto_accelerator.v:4224" *)
  wire _T_1499;
  (* src = "crypto_accelerator.v:4225" *)
  wire _T_1501;
  (* src = "crypto_accelerator.v:4226" *)
  wire _T_1503;
  (* src = "crypto_accelerator.v:4227" *)
  wire _T_1505;
  (* src = "crypto_accelerator.v:4228" *)
  wire _T_1507;
  (* src = "crypto_accelerator.v:4229" *)
  wire _T_1509;
  (* src = "crypto_accelerator.v:3558" *)
  wire _T_151;
  (* src = "crypto_accelerator.v:4230" *)
  wire _T_1511;
  (* src = "crypto_accelerator.v:4231" *)
  wire _T_1513;
  (* src = "crypto_accelerator.v:4232" *)
  wire _T_1515;
  (* src = "crypto_accelerator.v:4233" *)
  wire _T_1517;
  (* src = "crypto_accelerator.v:4234" *)
  wire _T_1519;
  (* src = "crypto_accelerator.v:4235" *)
  wire _T_1521;
  (* src = "crypto_accelerator.v:4236" *)
  wire _T_1523;
  (* src = "crypto_accelerator.v:4237" *)
  wire _T_1525;
  (* src = "crypto_accelerator.v:4238" *)
  wire _T_1527;
  (* src = "crypto_accelerator.v:4239" *)
  wire _T_1529;
  (* src = "crypto_accelerator.v:3559" *)
  wire _T_153;
  (* src = "crypto_accelerator.v:4240" *)
  wire _T_1531;
  (* src = "crypto_accelerator.v:4241" *)
  wire _T_1533;
  (* src = "crypto_accelerator.v:4242" *)
  wire _T_1535;
  (* src = "crypto_accelerator.v:4243" *)
  wire _T_1537;
  (* src = "crypto_accelerator.v:4244" *)
  wire _T_1539;
  (* src = "crypto_accelerator.v:4245" *)
  wire _T_1541;
  (* src = "crypto_accelerator.v:4246" *)
  wire _T_1543;
  (* src = "crypto_accelerator.v:4247" *)
  wire _T_1545;
  (* src = "crypto_accelerator.v:4248" *)
  wire _T_1547;
  (* src = "crypto_accelerator.v:4249" *)
  wire _T_1549;
  (* src = "crypto_accelerator.v:3560" *)
  wire _T_155;
  (* src = "crypto_accelerator.v:4250" *)
  wire _T_1551;
  (* src = "crypto_accelerator.v:4251" *)
  wire _T_1553;
  (* src = "crypto_accelerator.v:4252" *)
  wire _T_1555;
  (* src = "crypto_accelerator.v:4253" *)
  wire _T_1557;
  (* src = "crypto_accelerator.v:4254" *)
  wire _T_1559;
  (* src = "crypto_accelerator.v:4255" *)
  wire _T_1561;
  (* src = "crypto_accelerator.v:4256" *)
  wire _T_1563;
  (* src = "crypto_accelerator.v:4257" *)
  wire _T_1565;
  (* src = "crypto_accelerator.v:4258" *)
  wire _T_1567;
  (* src = "crypto_accelerator.v:4259" *)
  wire _T_1569;
  (* src = "crypto_accelerator.v:3561" *)
  wire _T_157;
  (* src = "crypto_accelerator.v:4260" *)
  wire _T_1571;
  (* src = "crypto_accelerator.v:4261" *)
  wire _T_1573;
  (* src = "crypto_accelerator.v:4262" *)
  wire _T_1575;
  (* src = "crypto_accelerator.v:4263" *)
  wire _T_1577;
  (* src = "crypto_accelerator.v:4264" *)
  wire _T_1579;
  (* src = "crypto_accelerator.v:4265" *)
  wire _T_1581;
  (* src = "crypto_accelerator.v:4266" *)
  wire _T_1583;
  (* src = "crypto_accelerator.v:4267" *)
  wire _T_1585;
  (* src = "crypto_accelerator.v:4268" *)
  wire _T_1587;
  (* src = "crypto_accelerator.v:4269" *)
  wire _T_1589;
  (* src = "crypto_accelerator.v:3562" *)
  wire _T_159;
  (* src = "crypto_accelerator.v:4270" *)
  wire _T_1591;
  (* src = "crypto_accelerator.v:4271" *)
  wire _T_1593;
  (* src = "crypto_accelerator.v:4272" *)
  wire _T_1595;
  (* src = "crypto_accelerator.v:4273" *)
  wire _T_1597;
  (* src = "crypto_accelerator.v:4274" *)
  wire _T_1599;
  (* src = "crypto_accelerator.v:4275" *)
  wire _T_1601;
  (* src = "crypto_accelerator.v:4276" *)
  wire _T_1603;
  (* src = "crypto_accelerator.v:4277" *)
  wire _T_1605;
  (* src = "crypto_accelerator.v:4278" *)
  wire _T_1607;
  (* src = "crypto_accelerator.v:4279" *)
  wire _T_1609;
  (* src = "crypto_accelerator.v:3563" *)
  wire _T_161;
  (* src = "crypto_accelerator.v:4280" *)
  wire _T_1611;
  (* src = "crypto_accelerator.v:4281" *)
  wire _T_1613;
  (* src = "crypto_accelerator.v:4282" *)
  wire _T_1615;
  (* src = "crypto_accelerator.v:4283" *)
  wire _T_1617;
  (* src = "crypto_accelerator.v:4284" *)
  wire _T_1619;
  (* src = "crypto_accelerator.v:4285" *)
  wire _T_1621;
  (* src = "crypto_accelerator.v:4286" *)
  wire _T_1623;
  (* src = "crypto_accelerator.v:4287" *)
  wire _T_1625;
  (* src = "crypto_accelerator.v:4288" *)
  wire _T_1627;
  (* src = "crypto_accelerator.v:4289" *)
  wire _T_1629;
  (* src = "crypto_accelerator.v:3564" *)
  wire _T_163;
  (* src = "crypto_accelerator.v:4290" *)
  wire _T_1631;
  (* src = "crypto_accelerator.v:4291" *)
  wire _T_1633;
  (* src = "crypto_accelerator.v:4292" *)
  wire _T_1635;
  (* src = "crypto_accelerator.v:4293" *)
  wire _T_1637;
  (* src = "crypto_accelerator.v:4294" *)
  wire _T_1639;
  (* src = "crypto_accelerator.v:4295" *)
  wire _T_1641;
  (* src = "crypto_accelerator.v:4296" *)
  wire _T_1643;
  (* src = "crypto_accelerator.v:4297" *)
  wire _T_1645;
  (* src = "crypto_accelerator.v:4298" *)
  wire _T_1647;
  (* src = "crypto_accelerator.v:4299" *)
  wire _T_1649;
  (* src = "crypto_accelerator.v:3565" *)
  wire _T_165;
  (* src = "crypto_accelerator.v:4300" *)
  wire _T_1651;
  (* src = "crypto_accelerator.v:4301" *)
  wire _T_1653;
  (* src = "crypto_accelerator.v:4302" *)
  wire _T_1655;
  (* src = "crypto_accelerator.v:4303" *)
  wire _T_1657;
  (* src = "crypto_accelerator.v:4304" *)
  wire _T_1659;
  (* src = "crypto_accelerator.v:4305" *)
  wire _T_1661;
  (* src = "crypto_accelerator.v:4306" *)
  wire _T_1663;
  (* src = "crypto_accelerator.v:4307" *)
  wire _T_1665;
  (* src = "crypto_accelerator.v:4308" *)
  wire _T_1667;
  (* src = "crypto_accelerator.v:4309" *)
  wire _T_1669;
  (* src = "crypto_accelerator.v:3566" *)
  wire _T_167;
  (* src = "crypto_accelerator.v:4310" *)
  wire _T_1671;
  (* src = "crypto_accelerator.v:4311" *)
  wire _T_1673;
  (* src = "crypto_accelerator.v:4312" *)
  wire _T_1675;
  (* src = "crypto_accelerator.v:4313" *)
  wire _T_1677;
  (* src = "crypto_accelerator.v:4314" *)
  wire _T_1679;
  (* src = "crypto_accelerator.v:4315" *)
  wire _T_1681;
  (* src = "crypto_accelerator.v:4316" *)
  wire _T_1683;
  (* src = "crypto_accelerator.v:4317" *)
  wire _T_1684;
  (* src = "crypto_accelerator.v:4318" *)
  wire _T_1685;
  (* src = "crypto_accelerator.v:4319" *)
  wire _T_1686;
  (* src = "crypto_accelerator.v:4320" *)
  wire _T_1687;
  (* src = "crypto_accelerator.v:4321" *)
  wire _T_1688;
  (* src = "crypto_accelerator.v:4322" *)
  wire _T_1689;
  (* src = "crypto_accelerator.v:3567" *)
  wire _T_169;
  (* src = "crypto_accelerator.v:4323" *)
  wire _T_1690;
  (* src = "crypto_accelerator.v:4324" *)
  wire _T_1691;
  (* src = "crypto_accelerator.v:3497" *)
  wire [63:0] _T_17;
  (* src = "crypto_accelerator.v:3568" *)
  wire _T_171;
  (* src = "crypto_accelerator.v:4326" *)
  wire _T_1716;
  (* src = "crypto_accelerator.v:4327" *)
  wire _T_1718;
  (* src = "crypto_accelerator.v:4328" *)
  wire _T_1719;
  (* src = "crypto_accelerator.v:4329" *)
  wire _T_1721;
  (* src = "crypto_accelerator.v:4330" *)
  wire _T_1722;
  (* src = "crypto_accelerator.v:4331" *)
  wire _T_1724;
  (* src = "crypto_accelerator.v:4332" *)
  wire _T_1726;
  (* src = "crypto_accelerator.v:4333" *)
  wire _T_1727;
  (* src = "crypto_accelerator.v:4334" *)
  wire _T_1729;
  (* src = "crypto_accelerator.v:3569" *)
  wire _T_173;
  (* src = "crypto_accelerator.v:4335" *)
  wire _T_1731;
  (* src = "crypto_accelerator.v:4336" *)
  wire _T_1732;
  (* src = "crypto_accelerator.v:4337" *)
  wire _T_1734;
  (* src = "crypto_accelerator.v:4338" *)
  wire _T_1736;
  (* src = "crypto_accelerator.v:4339" *)
  wire _T_1737;
  (* src = "crypto_accelerator.v:4340" *)
  wire _T_1739;
  (* src = "crypto_accelerator.v:4341" *)
  wire _T_1741;
  (* src = "crypto_accelerator.v:4342" *)
  wire _T_1743;
  (* src = "crypto_accelerator.v:4343" *)
  wire _T_1745;
  (* src = "crypto_accelerator.v:4344" *)
  wire _T_1746;
  (* src = "crypto_accelerator.v:4345" *)
  wire _T_1748;
  (* src = "crypto_accelerator.v:3570" *)
  wire _T_175;
  (* src = "crypto_accelerator.v:4346" *)
  wire _T_1750;
  (* src = "crypto_accelerator.v:4347" *)
  wire _T_1751;
  (* src = "crypto_accelerator.v:4348" *)
  wire _T_1753;
  (* src = "crypto_accelerator.v:4349" *)
  wire _T_1755;
  (* src = "crypto_accelerator.v:4350" *)
  wire _T_1757;
  (* src = "crypto_accelerator.v:4351" *)
  wire _T_1758;
  (* src = "crypto_accelerator.v:4352" *)
  wire _T_1760;
  (* src = "crypto_accelerator.v:4353" *)
  wire _T_1761;
  (* src = "crypto_accelerator.v:4354" *)
  wire _T_1763;
  (* src = "crypto_accelerator.v:4355" *)
  wire _T_1764;
  (* src = "crypto_accelerator.v:4356" *)
  wire _T_1766;
  (* src = "crypto_accelerator.v:4357" *)
  wire _T_1768;
  (* src = "crypto_accelerator.v:3571" *)
  wire _T_177;
  (* src = "crypto_accelerator.v:4358" *)
  wire _T_1770;
  (* src = "crypto_accelerator.v:4359" *)
  wire _T_1772;
  (* src = "crypto_accelerator.v:4360" *)
  wire _T_1774;
  (* src = "crypto_accelerator.v:4361" *)
  wire _T_1776;
  (* src = "crypto_accelerator.v:4362" *)
  wire _T_1778;
  (* src = "crypto_accelerator.v:4363" *)
  wire _T_1780;
  (* src = "crypto_accelerator.v:4364" *)
  wire _T_1782;
  (* src = "crypto_accelerator.v:4365" *)
  wire _T_1784;
  (* src = "crypto_accelerator.v:4366" *)
  wire _T_1786;
  (* src = "crypto_accelerator.v:4367" *)
  wire _T_1788;
  (* src = "crypto_accelerator.v:3572" *)
  wire _T_179;
  (* src = "crypto_accelerator.v:4368" *)
  wire _T_1790;
  (* src = "crypto_accelerator.v:4369" *)
  wire _T_1792;
  (* src = "crypto_accelerator.v:4370" *)
  wire _T_1794;
  (* src = "crypto_accelerator.v:4371" *)
  wire _T_1796;
  (* src = "crypto_accelerator.v:4372" *)
  wire _T_1798;
  (* src = "crypto_accelerator.v:4373" *)
  wire _T_1800;
  (* src = "crypto_accelerator.v:4374" *)
  wire _T_1802;
  (* src = "crypto_accelerator.v:4375" *)
  wire _T_1804;
  (* src = "crypto_accelerator.v:4376" *)
  wire _T_1806;
  (* src = "crypto_accelerator.v:4377" *)
  wire _T_1808;
  (* src = "crypto_accelerator.v:3573" *)
  wire _T_181;
  (* src = "crypto_accelerator.v:4378" *)
  wire _T_1810;
  (* src = "crypto_accelerator.v:4379" *)
  wire _T_1812;
  (* src = "crypto_accelerator.v:4380" *)
  wire _T_1814;
  (* src = "crypto_accelerator.v:4381" *)
  wire _T_1816;
  (* src = "crypto_accelerator.v:4382" *)
  wire _T_1818;
  (* src = "crypto_accelerator.v:4383" *)
  wire _T_1820;
  (* src = "crypto_accelerator.v:4384" *)
  wire _T_1822;
  (* src = "crypto_accelerator.v:4385" *)
  wire _T_1824;
  (* src = "crypto_accelerator.v:4386" *)
  wire _T_1826;
  (* src = "crypto_accelerator.v:4387" *)
  wire _T_1828;
  (* src = "crypto_accelerator.v:3574" *)
  wire _T_183;
  (* src = "crypto_accelerator.v:4388" *)
  wire _T_1830;
  (* src = "crypto_accelerator.v:4389" *)
  wire _T_1832;
  (* src = "crypto_accelerator.v:4390" *)
  wire _T_1834;
  (* src = "crypto_accelerator.v:4391" *)
  wire _T_1836;
  (* src = "crypto_accelerator.v:4392" *)
  wire _T_1838;
  (* src = "crypto_accelerator.v:4393" *)
  wire _T_1840;
  (* src = "crypto_accelerator.v:4394" *)
  wire _T_1842;
  (* src = "crypto_accelerator.v:4395" *)
  wire _T_1844;
  (* src = "crypto_accelerator.v:4396" *)
  wire _T_1846;
  (* src = "crypto_accelerator.v:4397" *)
  wire _T_1848;
  (* src = "crypto_accelerator.v:3575" *)
  wire _T_185;
  (* src = "crypto_accelerator.v:4398" *)
  wire _T_1850;
  (* src = "crypto_accelerator.v:4399" *)
  wire _T_1852;
  (* src = "crypto_accelerator.v:4400" *)
  wire _T_1854;
  (* src = "crypto_accelerator.v:4401" *)
  wire _T_1856;
  (* src = "crypto_accelerator.v:4402" *)
  wire _T_1858;
  (* src = "crypto_accelerator.v:4403" *)
  wire _T_1860;
  (* src = "crypto_accelerator.v:4404" *)
  wire _T_1862;
  (* src = "crypto_accelerator.v:4405" *)
  wire _T_1864;
  (* src = "crypto_accelerator.v:4406" *)
  wire _T_1866;
  (* src = "crypto_accelerator.v:4407" *)
  wire _T_1868;
  (* src = "crypto_accelerator.v:3576" *)
  wire _T_187;
  (* src = "crypto_accelerator.v:4408" *)
  wire _T_1870;
  (* src = "crypto_accelerator.v:4409" *)
  wire _T_1872;
  (* src = "crypto_accelerator.v:4410" *)
  wire _T_1874;
  (* src = "crypto_accelerator.v:4411" *)
  wire _T_1876;
  (* src = "crypto_accelerator.v:4412" *)
  wire _T_1878;
  (* src = "crypto_accelerator.v:4413" *)
  wire _T_1880;
  (* src = "crypto_accelerator.v:4414" *)
  wire _T_1882;
  (* src = "crypto_accelerator.v:4415" *)
  wire _T_1884;
  (* src = "crypto_accelerator.v:4416" *)
  wire _T_1886;
  (* src = "crypto_accelerator.v:4417" *)
  wire _T_1888;
  (* src = "crypto_accelerator.v:3577" *)
  wire _T_189;
  (* src = "crypto_accelerator.v:4418" *)
  wire _T_1890;
  (* src = "crypto_accelerator.v:4419" *)
  wire _T_1892;
  (* src = "crypto_accelerator.v:4420" *)
  wire _T_1894;
  (* src = "crypto_accelerator.v:4421" *)
  wire _T_1896;
  (* src = "crypto_accelerator.v:4422" *)
  wire _T_1898;
  (* src = "crypto_accelerator.v:4423" *)
  wire _T_1900;
  (* src = "crypto_accelerator.v:4424" *)
  wire _T_1902;
  (* src = "crypto_accelerator.v:4425" *)
  wire _T_1904;
  (* src = "crypto_accelerator.v:4426" *)
  wire _T_1906;
  (* src = "crypto_accelerator.v:4427" *)
  wire _T_1908;
  (* src = "crypto_accelerator.v:3578" *)
  wire _T_191;
  (* src = "crypto_accelerator.v:4428" *)
  wire _T_1910;
  (* src = "crypto_accelerator.v:4429" *)
  wire _T_1912;
  (* src = "crypto_accelerator.v:4430" *)
  wire _T_1914;
  (* src = "crypto_accelerator.v:4431" *)
  wire _T_1916;
  (* src = "crypto_accelerator.v:4432" *)
  wire _T_1918;
  (* src = "crypto_accelerator.v:4433" *)
  wire _T_1920;
  (* src = "crypto_accelerator.v:4434" *)
  wire _T_1922;
  (* src = "crypto_accelerator.v:4435" *)
  wire _T_1924;
  (* src = "crypto_accelerator.v:4436" *)
  wire _T_1926;
  (* src = "crypto_accelerator.v:4437" *)
  wire _T_1928;
  (* src = "crypto_accelerator.v:3579" *)
  wire _T_193;
  (* src = "crypto_accelerator.v:4438" *)
  wire _T_1930;
  (* src = "crypto_accelerator.v:4439" *)
  wire _T_1932;
  (* src = "crypto_accelerator.v:4440" *)
  wire _T_1934;
  (* src = "crypto_accelerator.v:4441" *)
  wire _T_1936;
  (* src = "crypto_accelerator.v:4442" *)
  wire _T_1938;
  (* src = "crypto_accelerator.v:4443" *)
  wire _T_1940;
  (* src = "crypto_accelerator.v:4444" *)
  wire _T_1942;
  (* src = "crypto_accelerator.v:4445" *)
  wire _T_1944;
  (* src = "crypto_accelerator.v:4446" *)
  wire _T_1946;
  (* src = "crypto_accelerator.v:4447" *)
  wire _T_1948;
  (* src = "crypto_accelerator.v:3580" *)
  wire _T_195;
  (* src = "crypto_accelerator.v:4448" *)
  wire _T_1950;
  (* src = "crypto_accelerator.v:4449" *)
  wire _T_1952;
  (* src = "crypto_accelerator.v:4450" *)
  wire _T_1954;
  (* src = "crypto_accelerator.v:4451" *)
  wire _T_1956;
  (* src = "crypto_accelerator.v:4452" *)
  wire _T_1958;
  (* src = "crypto_accelerator.v:4453" *)
  wire _T_1960;
  (* src = "crypto_accelerator.v:4454" *)
  wire _T_1962;
  (* src = "crypto_accelerator.v:4455" *)
  wire _T_1963;
  (* src = "crypto_accelerator.v:4456" *)
  wire _T_1964;
  (* src = "crypto_accelerator.v:4457" *)
  wire _T_1965;
  (* src = "crypto_accelerator.v:4458" *)
  wire _T_1966;
  (* src = "crypto_accelerator.v:4459" *)
  wire _T_1967;
  (* src = "crypto_accelerator.v:4460" *)
  wire _T_1968;
  (* src = "crypto_accelerator.v:4461" *)
  wire _T_1969;
  (* src = "crypto_accelerator.v:3581" *)
  wire _T_197;
  (* src = "crypto_accelerator.v:4462" *)
  wire _T_1970;
  (* src = "crypto_accelerator.v:3582" *)
  wire _T_199;
  (* src = "crypto_accelerator.v:4464" *)
  wire _T_1995;
  (* src = "crypto_accelerator.v:4465" *)
  wire _T_1997;
  (* src = "crypto_accelerator.v:4466" *)
  wire _T_1998;
  (* src = "crypto_accelerator.v:4467" *)
  wire _T_2000;
  (* src = "crypto_accelerator.v:4468" *)
  wire _T_2001;
  (* src = "crypto_accelerator.v:4469" *)
  wire _T_2003;
  (* src = "crypto_accelerator.v:4470" *)
  wire _T_2005;
  (* src = "crypto_accelerator.v:4471" *)
  wire _T_2006;
  (* src = "crypto_accelerator.v:4472" *)
  wire _T_2008;
  (* src = "crypto_accelerator.v:3583" *)
  wire _T_201;
  (* src = "crypto_accelerator.v:4473" *)
  wire _T_2010;
  (* src = "crypto_accelerator.v:4474" *)
  wire _T_2011;
  (* src = "crypto_accelerator.v:4475" *)
  wire _T_2013;
  (* src = "crypto_accelerator.v:4476" *)
  wire _T_2015;
  (* src = "crypto_accelerator.v:4477" *)
  wire _T_2016;
  (* src = "crypto_accelerator.v:4478" *)
  wire _T_2018;
  (* src = "crypto_accelerator.v:4479" *)
  wire _T_2020;
  (* src = "crypto_accelerator.v:4480" *)
  wire _T_2022;
  (* src = "crypto_accelerator.v:4481" *)
  wire _T_2024;
  (* src = "crypto_accelerator.v:4482" *)
  wire _T_2025;
  (* src = "crypto_accelerator.v:4483" *)
  wire _T_2027;
  (* src = "crypto_accelerator.v:4484" *)
  wire _T_2029;
  (* src = "crypto_accelerator.v:3584" *)
  wire _T_203;
  (* src = "crypto_accelerator.v:4485" *)
  wire _T_2030;
  (* src = "crypto_accelerator.v:4486" *)
  wire _T_2032;
  (* src = "crypto_accelerator.v:4487" *)
  wire _T_2034;
  (* src = "crypto_accelerator.v:4488" *)
  wire _T_2036;
  (* src = "crypto_accelerator.v:4489" *)
  wire _T_2037;
  (* src = "crypto_accelerator.v:4490" *)
  wire _T_2039;
  (* src = "crypto_accelerator.v:4491" *)
  wire _T_2040;
  (* src = "crypto_accelerator.v:4492" *)
  wire _T_2042;
  (* src = "crypto_accelerator.v:4493" *)
  wire _T_2043;
  (* src = "crypto_accelerator.v:4494" *)
  wire _T_2045;
  (* src = "crypto_accelerator.v:4495" *)
  wire _T_2047;
  (* src = "crypto_accelerator.v:4496" *)
  wire _T_2049;
  (* src = "crypto_accelerator.v:3585" *)
  wire _T_205;
  (* src = "crypto_accelerator.v:4497" *)
  wire _T_2051;
  (* src = "crypto_accelerator.v:4498" *)
  wire _T_2053;
  (* src = "crypto_accelerator.v:4499" *)
  wire _T_2055;
  (* src = "crypto_accelerator.v:4500" *)
  wire _T_2057;
  (* src = "crypto_accelerator.v:4501" *)
  wire _T_2059;
  (* src = "crypto_accelerator.v:4502" *)
  wire _T_2061;
  (* src = "crypto_accelerator.v:4503" *)
  wire _T_2063;
  (* src = "crypto_accelerator.v:4504" *)
  wire _T_2065;
  (* src = "crypto_accelerator.v:4505" *)
  wire _T_2067;
  (* src = "crypto_accelerator.v:4506" *)
  wire _T_2069;
  (* src = "crypto_accelerator.v:3586" *)
  wire _T_207;
  (* src = "crypto_accelerator.v:4507" *)
  wire _T_2071;
  (* src = "crypto_accelerator.v:4508" *)
  wire _T_2073;
  (* src = "crypto_accelerator.v:4509" *)
  wire _T_2075;
  (* src = "crypto_accelerator.v:4510" *)
  wire _T_2077;
  (* src = "crypto_accelerator.v:4511" *)
  wire _T_2079;
  (* src = "crypto_accelerator.v:4512" *)
  wire _T_2081;
  (* src = "crypto_accelerator.v:4513" *)
  wire _T_2083;
  (* src = "crypto_accelerator.v:4514" *)
  wire _T_2085;
  (* src = "crypto_accelerator.v:4515" *)
  wire _T_2087;
  (* src = "crypto_accelerator.v:4516" *)
  wire _T_2089;
  (* src = "crypto_accelerator.v:3587" *)
  wire _T_209;
  (* src = "crypto_accelerator.v:4517" *)
  wire _T_2091;
  (* src = "crypto_accelerator.v:4518" *)
  wire _T_2093;
  (* src = "crypto_accelerator.v:4519" *)
  wire _T_2095;
  (* src = "crypto_accelerator.v:4520" *)
  wire _T_2097;
  (* src = "crypto_accelerator.v:4521" *)
  wire _T_2099;
  (* src = "crypto_accelerator.v:4522" *)
  wire _T_2101;
  (* src = "crypto_accelerator.v:4523" *)
  wire _T_2103;
  (* src = "crypto_accelerator.v:4524" *)
  wire _T_2105;
  (* src = "crypto_accelerator.v:4525" *)
  wire _T_2107;
  (* src = "crypto_accelerator.v:4526" *)
  wire _T_2109;
  (* src = "crypto_accelerator.v:3588" *)
  wire _T_211;
  (* src = "crypto_accelerator.v:4527" *)
  wire _T_2111;
  (* src = "crypto_accelerator.v:4528" *)
  wire _T_2113;
  (* src = "crypto_accelerator.v:4529" *)
  wire _T_2115;
  (* src = "crypto_accelerator.v:4530" *)
  wire _T_2117;
  (* src = "crypto_accelerator.v:4531" *)
  wire _T_2119;
  (* src = "crypto_accelerator.v:4532" *)
  wire _T_2121;
  (* src = "crypto_accelerator.v:4533" *)
  wire _T_2123;
  (* src = "crypto_accelerator.v:4534" *)
  wire _T_2125;
  (* src = "crypto_accelerator.v:4535" *)
  wire _T_2127;
  (* src = "crypto_accelerator.v:4536" *)
  wire _T_2129;
  (* src = "crypto_accelerator.v:3589" *)
  wire _T_213;
  (* src = "crypto_accelerator.v:4537" *)
  wire _T_2131;
  (* src = "crypto_accelerator.v:4538" *)
  wire _T_2133;
  (* src = "crypto_accelerator.v:4539" *)
  wire _T_2135;
  (* src = "crypto_accelerator.v:4540" *)
  wire _T_2137;
  (* src = "crypto_accelerator.v:4541" *)
  wire _T_2139;
  (* src = "crypto_accelerator.v:4542" *)
  wire _T_2141;
  (* src = "crypto_accelerator.v:4543" *)
  wire _T_2143;
  (* src = "crypto_accelerator.v:4544" *)
  wire _T_2145;
  (* src = "crypto_accelerator.v:4545" *)
  wire _T_2147;
  (* src = "crypto_accelerator.v:4546" *)
  wire _T_2149;
  (* src = "crypto_accelerator.v:3590" *)
  wire _T_215;
  (* src = "crypto_accelerator.v:4547" *)
  wire _T_2151;
  (* src = "crypto_accelerator.v:4548" *)
  wire _T_2153;
  (* src = "crypto_accelerator.v:4549" *)
  wire _T_2155;
  (* src = "crypto_accelerator.v:4550" *)
  wire _T_2157;
  (* src = "crypto_accelerator.v:4551" *)
  wire _T_2159;
  (* src = "crypto_accelerator.v:4552" *)
  wire _T_2161;
  (* src = "crypto_accelerator.v:4553" *)
  wire _T_2163;
  (* src = "crypto_accelerator.v:4554" *)
  wire _T_2165;
  (* src = "crypto_accelerator.v:4555" *)
  wire _T_2167;
  (* src = "crypto_accelerator.v:4556" *)
  wire _T_2169;
  (* src = "crypto_accelerator.v:3591" *)
  wire _T_217;
  (* src = "crypto_accelerator.v:4557" *)
  wire _T_2171;
  (* src = "crypto_accelerator.v:4558" *)
  wire _T_2173;
  (* src = "crypto_accelerator.v:4559" *)
  wire _T_2175;
  (* src = "crypto_accelerator.v:4560" *)
  wire _T_2177;
  (* src = "crypto_accelerator.v:4561" *)
  wire _T_2179;
  (* src = "crypto_accelerator.v:4562" *)
  wire _T_2181;
  (* src = "crypto_accelerator.v:4563" *)
  wire _T_2183;
  (* src = "crypto_accelerator.v:4564" *)
  wire _T_2185;
  (* src = "crypto_accelerator.v:4565" *)
  wire _T_2187;
  (* src = "crypto_accelerator.v:4566" *)
  wire _T_2189;
  (* src = "crypto_accelerator.v:3592" *)
  wire _T_219;
  (* src = "crypto_accelerator.v:4567" *)
  wire _T_2191;
  (* src = "crypto_accelerator.v:4568" *)
  wire _T_2193;
  (* src = "crypto_accelerator.v:4569" *)
  wire _T_2195;
  (* src = "crypto_accelerator.v:4570" *)
  wire _T_2197;
  (* src = "crypto_accelerator.v:4571" *)
  wire _T_2199;
  (* src = "crypto_accelerator.v:4572" *)
  wire _T_2201;
  (* src = "crypto_accelerator.v:4573" *)
  wire _T_2203;
  (* src = "crypto_accelerator.v:4574" *)
  wire _T_2205;
  (* src = "crypto_accelerator.v:4575" *)
  wire _T_2207;
  (* src = "crypto_accelerator.v:4576" *)
  wire _T_2209;
  (* src = "crypto_accelerator.v:3593" *)
  wire _T_221;
  (* src = "crypto_accelerator.v:4577" *)
  wire _T_2211;
  (* src = "crypto_accelerator.v:4578" *)
  wire _T_2213;
  (* src = "crypto_accelerator.v:4579" *)
  wire _T_2215;
  (* src = "crypto_accelerator.v:4580" *)
  wire _T_2217;
  (* src = "crypto_accelerator.v:4581" *)
  wire _T_2219;
  (* src = "crypto_accelerator.v:4582" *)
  wire _T_2221;
  (* src = "crypto_accelerator.v:4583" *)
  wire _T_2223;
  (* src = "crypto_accelerator.v:4584" *)
  wire _T_2225;
  (* src = "crypto_accelerator.v:4585" *)
  wire _T_2227;
  (* src = "crypto_accelerator.v:4586" *)
  wire _T_2229;
  (* src = "crypto_accelerator.v:3594" *)
  wire _T_223;
  (* src = "crypto_accelerator.v:4587" *)
  wire _T_2231;
  (* src = "crypto_accelerator.v:4588" *)
  wire _T_2233;
  (* src = "crypto_accelerator.v:4589" *)
  wire _T_2235;
  (* src = "crypto_accelerator.v:4590" *)
  wire _T_2237;
  (* src = "crypto_accelerator.v:4591" *)
  wire _T_2239;
  (* src = "crypto_accelerator.v:4592" *)
  wire _T_2241;
  (* src = "crypto_accelerator.v:4593" *)
  wire _T_2242;
  (* src = "crypto_accelerator.v:4594" *)
  wire _T_2243;
  (* src = "crypto_accelerator.v:4595" *)
  wire _T_2244;
  (* src = "crypto_accelerator.v:4596" *)
  wire _T_2245;
  (* src = "crypto_accelerator.v:4597" *)
  wire _T_2246;
  (* src = "crypto_accelerator.v:4598" *)
  wire _T_2247;
  (* src = "crypto_accelerator.v:4599" *)
  wire _T_2248;
  (* src = "crypto_accelerator.v:4600" *)
  wire _T_2249;
  (* src = "crypto_accelerator.v:3595" *)
  wire _T_225;
  (* src = "crypto_accelerator.v:3596" *)
  wire _T_227;
  (* src = "crypto_accelerator.v:4602" *)
  wire _T_2275;
  (* src = "crypto_accelerator.v:4603" *)
  wire _T_2277;
  (* src = "crypto_accelerator.v:4604" *)
  wire _T_2278;
  (* src = "crypto_accelerator.v:4605" *)
  wire _T_2280;
  (* src = "crypto_accelerator.v:4606" *)
  wire _T_2281;
  (* src = "crypto_accelerator.v:4607" *)
  wire _T_2283;
  (* src = "crypto_accelerator.v:4608" *)
  wire _T_2285;
  (* src = "crypto_accelerator.v:4609" *)
  wire _T_2286;
  (* src = "crypto_accelerator.v:4610" *)
  wire _T_2288;
  (* src = "crypto_accelerator.v:3597" *)
  wire _T_229;
  (* src = "crypto_accelerator.v:4611" *)
  wire _T_2290;
  (* src = "crypto_accelerator.v:4612" *)
  wire _T_2291;
  (* src = "crypto_accelerator.v:4613" *)
  wire _T_2293;
  (* src = "crypto_accelerator.v:4614" *)
  wire _T_2295;
  (* src = "crypto_accelerator.v:4615" *)
  wire _T_2296;
  (* src = "crypto_accelerator.v:4616" *)
  wire _T_2298;
  (* src = "crypto_accelerator.v:4617" *)
  wire _T_2300;
  (* src = "crypto_accelerator.v:4618" *)
  wire _T_2302;
  (* src = "crypto_accelerator.v:4619" *)
  wire _T_2304;
  (* src = "crypto_accelerator.v:4620" *)
  wire _T_2305;
  (* src = "crypto_accelerator.v:4621" *)
  wire _T_2307;
  (* src = "crypto_accelerator.v:4622" *)
  wire _T_2309;
  (* src = "crypto_accelerator.v:3598" *)
  wire _T_231;
  (* src = "crypto_accelerator.v:4623" *)
  wire _T_2310;
  (* src = "crypto_accelerator.v:4624" *)
  wire _T_2312;
  (* src = "crypto_accelerator.v:4625" *)
  wire _T_2314;
  (* src = "crypto_accelerator.v:4626" *)
  wire _T_2316;
  (* src = "crypto_accelerator.v:4627" *)
  wire _T_2317;
  (* src = "crypto_accelerator.v:4628" *)
  wire _T_2319;
  (* src = "crypto_accelerator.v:4629" *)
  wire _T_2320;
  (* src = "crypto_accelerator.v:4630" *)
  wire _T_2322;
  (* src = "crypto_accelerator.v:4631" *)
  wire _T_2323;
  (* src = "crypto_accelerator.v:4632" *)
  wire _T_2325;
  (* src = "crypto_accelerator.v:4633" *)
  wire _T_2327;
  (* src = "crypto_accelerator.v:4634" *)
  wire _T_2329;
  (* src = "crypto_accelerator.v:3599" *)
  wire _T_233;
  (* src = "crypto_accelerator.v:4635" *)
  wire _T_2331;
  (* src = "crypto_accelerator.v:4636" *)
  wire _T_2333;
  (* src = "crypto_accelerator.v:4637" *)
  wire _T_2335;
  (* src = "crypto_accelerator.v:4638" *)
  wire _T_2337;
  (* src = "crypto_accelerator.v:4639" *)
  wire _T_2339;
  (* src = "crypto_accelerator.v:4640" *)
  wire _T_2341;
  (* src = "crypto_accelerator.v:4641" *)
  wire _T_2343;
  (* src = "crypto_accelerator.v:4642" *)
  wire _T_2345;
  (* src = "crypto_accelerator.v:4643" *)
  wire _T_2347;
  (* src = "crypto_accelerator.v:4644" *)
  wire _T_2349;
  (* src = "crypto_accelerator.v:3600" *)
  wire _T_235;
  (* src = "crypto_accelerator.v:4645" *)
  wire _T_2351;
  (* src = "crypto_accelerator.v:4646" *)
  wire _T_2353;
  (* src = "crypto_accelerator.v:4647" *)
  wire _T_2355;
  (* src = "crypto_accelerator.v:4648" *)
  wire _T_2357;
  (* src = "crypto_accelerator.v:4649" *)
  wire _T_2359;
  (* src = "crypto_accelerator.v:4650" *)
  wire _T_2361;
  (* src = "crypto_accelerator.v:4651" *)
  wire _T_2363;
  (* src = "crypto_accelerator.v:4652" *)
  wire _T_2365;
  (* src = "crypto_accelerator.v:4653" *)
  wire _T_2367;
  (* src = "crypto_accelerator.v:4654" *)
  wire _T_2369;
  (* src = "crypto_accelerator.v:3601" *)
  wire _T_237;
  (* src = "crypto_accelerator.v:4655" *)
  wire _T_2371;
  (* src = "crypto_accelerator.v:4656" *)
  wire _T_2373;
  (* src = "crypto_accelerator.v:4657" *)
  wire _T_2375;
  (* src = "crypto_accelerator.v:4658" *)
  wire _T_2377;
  (* src = "crypto_accelerator.v:4659" *)
  wire _T_2379;
  (* src = "crypto_accelerator.v:4660" *)
  wire _T_2381;
  (* src = "crypto_accelerator.v:4661" *)
  wire _T_2383;
  (* src = "crypto_accelerator.v:4662" *)
  wire _T_2385;
  (* src = "crypto_accelerator.v:4663" *)
  wire _T_2387;
  (* src = "crypto_accelerator.v:4664" *)
  wire _T_2389;
  (* src = "crypto_accelerator.v:3602" *)
  wire _T_239;
  (* src = "crypto_accelerator.v:4665" *)
  wire _T_2391;
  (* src = "crypto_accelerator.v:4666" *)
  wire _T_2393;
  (* src = "crypto_accelerator.v:4667" *)
  wire _T_2395;
  (* src = "crypto_accelerator.v:4668" *)
  wire _T_2397;
  (* src = "crypto_accelerator.v:4669" *)
  wire _T_2399;
  (* src = "crypto_accelerator.v:4670" *)
  wire _T_2401;
  (* src = "crypto_accelerator.v:4671" *)
  wire _T_2403;
  (* src = "crypto_accelerator.v:4672" *)
  wire _T_2405;
  (* src = "crypto_accelerator.v:4673" *)
  wire _T_2407;
  (* src = "crypto_accelerator.v:4674" *)
  wire _T_2409;
  (* src = "crypto_accelerator.v:3603" *)
  wire _T_241;
  (* src = "crypto_accelerator.v:4675" *)
  wire _T_2411;
  (* src = "crypto_accelerator.v:4676" *)
  wire _T_2413;
  (* src = "crypto_accelerator.v:4677" *)
  wire _T_2415;
  (* src = "crypto_accelerator.v:4678" *)
  wire _T_2417;
  (* src = "crypto_accelerator.v:4679" *)
  wire _T_2419;
  (* src = "crypto_accelerator.v:4680" *)
  wire _T_2421;
  (* src = "crypto_accelerator.v:4681" *)
  wire _T_2423;
  (* src = "crypto_accelerator.v:4682" *)
  wire _T_2425;
  (* src = "crypto_accelerator.v:4683" *)
  wire _T_2427;
  (* src = "crypto_accelerator.v:4684" *)
  wire _T_2429;
  (* src = "crypto_accelerator.v:3604" *)
  wire _T_243;
  (* src = "crypto_accelerator.v:4685" *)
  wire _T_2431;
  (* src = "crypto_accelerator.v:4686" *)
  wire _T_2433;
  (* src = "crypto_accelerator.v:4687" *)
  wire _T_2435;
  (* src = "crypto_accelerator.v:4688" *)
  wire _T_2437;
  (* src = "crypto_accelerator.v:4689" *)
  wire _T_2439;
  (* src = "crypto_accelerator.v:4690" *)
  wire _T_2441;
  (* src = "crypto_accelerator.v:4691" *)
  wire _T_2443;
  (* src = "crypto_accelerator.v:4692" *)
  wire _T_2445;
  (* src = "crypto_accelerator.v:4693" *)
  wire _T_2447;
  (* src = "crypto_accelerator.v:4694" *)
  wire _T_2449;
  (* src = "crypto_accelerator.v:3605" *)
  wire _T_245;
  (* src = "crypto_accelerator.v:4695" *)
  wire _T_2451;
  (* src = "crypto_accelerator.v:4696" *)
  wire _T_2453;
  (* src = "crypto_accelerator.v:4697" *)
  wire _T_2455;
  (* src = "crypto_accelerator.v:4698" *)
  wire _T_2457;
  (* src = "crypto_accelerator.v:4699" *)
  wire _T_2459;
  (* src = "crypto_accelerator.v:4700" *)
  wire _T_2461;
  (* src = "crypto_accelerator.v:4701" *)
  wire _T_2463;
  (* src = "crypto_accelerator.v:4702" *)
  wire _T_2465;
  (* src = "crypto_accelerator.v:4703" *)
  wire _T_2467;
  (* src = "crypto_accelerator.v:4704" *)
  wire _T_2469;
  (* src = "crypto_accelerator.v:3606" *)
  wire _T_247;
  (* src = "crypto_accelerator.v:4705" *)
  wire _T_2471;
  (* src = "crypto_accelerator.v:4706" *)
  wire _T_2473;
  (* src = "crypto_accelerator.v:4707" *)
  wire _T_2475;
  (* src = "crypto_accelerator.v:4708" *)
  wire _T_2477;
  (* src = "crypto_accelerator.v:4709" *)
  wire _T_2479;
  (* src = "crypto_accelerator.v:4710" *)
  wire _T_2481;
  (* src = "crypto_accelerator.v:4711" *)
  wire _T_2483;
  (* src = "crypto_accelerator.v:4712" *)
  wire _T_2485;
  (* src = "crypto_accelerator.v:4713" *)
  wire _T_2487;
  (* src = "crypto_accelerator.v:4714" *)
  wire _T_2489;
  (* src = "crypto_accelerator.v:3607" *)
  wire _T_249;
  (* src = "crypto_accelerator.v:4715" *)
  wire _T_2491;
  (* src = "crypto_accelerator.v:4716" *)
  wire _T_2493;
  (* src = "crypto_accelerator.v:4717" *)
  wire _T_2495;
  (* src = "crypto_accelerator.v:4718" *)
  wire _T_2497;
  (* src = "crypto_accelerator.v:4719" *)
  wire _T_2499;
  (* src = "crypto_accelerator.v:4720" *)
  wire _T_2501;
  (* src = "crypto_accelerator.v:4721" *)
  wire _T_2503;
  (* src = "crypto_accelerator.v:4722" *)
  wire _T_2505;
  (* src = "crypto_accelerator.v:4723" *)
  wire _T_2507;
  (* src = "crypto_accelerator.v:4724" *)
  wire _T_2509;
  (* src = "crypto_accelerator.v:3608" *)
  wire _T_251;
  (* src = "crypto_accelerator.v:4725" *)
  wire _T_2511;
  (* src = "crypto_accelerator.v:4726" *)
  wire _T_2513;
  (* src = "crypto_accelerator.v:4727" *)
  wire _T_2515;
  (* src = "crypto_accelerator.v:4728" *)
  wire _T_2517;
  (* src = "crypto_accelerator.v:4729" *)
  wire _T_2519;
  (* src = "crypto_accelerator.v:4730" *)
  wire _T_2521;
  (* src = "crypto_accelerator.v:4731" *)
  wire _T_2522;
  (* src = "crypto_accelerator.v:4732" *)
  wire _T_2523;
  (* src = "crypto_accelerator.v:4733" *)
  wire _T_2524;
  (* src = "crypto_accelerator.v:4734" *)
  wire _T_2525;
  (* src = "crypto_accelerator.v:4735" *)
  wire _T_2526;
  (* src = "crypto_accelerator.v:4736" *)
  wire _T_2527;
  (* src = "crypto_accelerator.v:4737" *)
  wire _T_2528;
  (* src = "crypto_accelerator.v:4738" *)
  wire _T_2529;
  (* src = "crypto_accelerator.v:3609" *)
  wire _T_253;
  (* src = "crypto_accelerator.v:3610" *)
  wire _T_255;
  (* src = "crypto_accelerator.v:4740" *)
  wire _T_2554;
  (* src = "crypto_accelerator.v:4741" *)
  wire _T_2556;
  (* src = "crypto_accelerator.v:4742" *)
  wire _T_2557;
  (* src = "crypto_accelerator.v:4743" *)
  wire _T_2559;
  (* src = "crypto_accelerator.v:4744" *)
  wire _T_2560;
  (* src = "crypto_accelerator.v:4745" *)
  wire _T_2562;
  (* src = "crypto_accelerator.v:4746" *)
  wire _T_2564;
  (* src = "crypto_accelerator.v:4747" *)
  wire _T_2565;
  (* src = "crypto_accelerator.v:4748" *)
  wire _T_2567;
  (* src = "crypto_accelerator.v:4749" *)
  wire _T_2569;
  (* src = "crypto_accelerator.v:3611" *)
  wire _T_257;
  (* src = "crypto_accelerator.v:4750" *)
  wire _T_2570;
  (* src = "crypto_accelerator.v:4751" *)
  wire _T_2572;
  (* src = "crypto_accelerator.v:4752" *)
  wire _T_2574;
  (* src = "crypto_accelerator.v:4753" *)
  wire _T_2575;
  (* src = "crypto_accelerator.v:4754" *)
  wire _T_2577;
  (* src = "crypto_accelerator.v:4755" *)
  wire _T_2579;
  (* src = "crypto_accelerator.v:4756" *)
  wire _T_2581;
  (* src = "crypto_accelerator.v:4757" *)
  wire _T_2583;
  (* src = "crypto_accelerator.v:4758" *)
  wire _T_2584;
  (* src = "crypto_accelerator.v:4759" *)
  wire _T_2586;
  (* src = "crypto_accelerator.v:4760" *)
  wire _T_2588;
  (* src = "crypto_accelerator.v:4761" *)
  wire _T_2589;
  (* src = "crypto_accelerator.v:3612" *)
  wire _T_259;
  (* src = "crypto_accelerator.v:4762" *)
  wire _T_2591;
  (* src = "crypto_accelerator.v:4763" *)
  wire _T_2593;
  (* src = "crypto_accelerator.v:4764" *)
  wire _T_2595;
  (* src = "crypto_accelerator.v:4765" *)
  wire _T_2596;
  (* src = "crypto_accelerator.v:4766" *)
  wire _T_2598;
  (* src = "crypto_accelerator.v:4767" *)
  wire _T_2599;
  (* src = "crypto_accelerator.v:4768" *)
  wire _T_2601;
  (* src = "crypto_accelerator.v:4769" *)
  wire _T_2602;
  (* src = "crypto_accelerator.v:4770" *)
  wire _T_2604;
  (* src = "crypto_accelerator.v:4771" *)
  wire _T_2606;
  (* src = "crypto_accelerator.v:4772" *)
  wire _T_2608;
  (* src = "crypto_accelerator.v:3613" *)
  wire _T_261;
  (* src = "crypto_accelerator.v:4773" *)
  wire _T_2610;
  (* src = "crypto_accelerator.v:4774" *)
  wire _T_2612;
  (* src = "crypto_accelerator.v:4775" *)
  wire _T_2614;
  (* src = "crypto_accelerator.v:4776" *)
  wire _T_2616;
  (* src = "crypto_accelerator.v:4777" *)
  wire _T_2618;
  (* src = "crypto_accelerator.v:4778" *)
  wire _T_2620;
  (* src = "crypto_accelerator.v:4779" *)
  wire _T_2622;
  (* src = "crypto_accelerator.v:4780" *)
  wire _T_2624;
  (* src = "crypto_accelerator.v:4781" *)
  wire _T_2626;
  (* src = "crypto_accelerator.v:4782" *)
  wire _T_2628;
  (* src = "crypto_accelerator.v:3614" *)
  wire _T_263;
  (* src = "crypto_accelerator.v:4783" *)
  wire _T_2630;
  (* src = "crypto_accelerator.v:4784" *)
  wire _T_2632;
  (* src = "crypto_accelerator.v:4785" *)
  wire _T_2634;
  (* src = "crypto_accelerator.v:4786" *)
  wire _T_2636;
  (* src = "crypto_accelerator.v:4787" *)
  wire _T_2638;
  (* src = "crypto_accelerator.v:4788" *)
  wire _T_2640;
  (* src = "crypto_accelerator.v:4789" *)
  wire _T_2642;
  (* src = "crypto_accelerator.v:4790" *)
  wire _T_2644;
  (* src = "crypto_accelerator.v:4791" *)
  wire _T_2646;
  (* src = "crypto_accelerator.v:4792" *)
  wire _T_2648;
  (* src = "crypto_accelerator.v:3615" *)
  wire _T_265;
  (* src = "crypto_accelerator.v:4793" *)
  wire _T_2650;
  (* src = "crypto_accelerator.v:4794" *)
  wire _T_2652;
  (* src = "crypto_accelerator.v:4795" *)
  wire _T_2654;
  (* src = "crypto_accelerator.v:4796" *)
  wire _T_2656;
  (* src = "crypto_accelerator.v:4797" *)
  wire _T_2658;
  (* src = "crypto_accelerator.v:4798" *)
  wire _T_2660;
  (* src = "crypto_accelerator.v:4799" *)
  wire _T_2662;
  (* src = "crypto_accelerator.v:4800" *)
  wire _T_2664;
  (* src = "crypto_accelerator.v:4801" *)
  wire _T_2666;
  (* src = "crypto_accelerator.v:4802" *)
  wire _T_2668;
  (* src = "crypto_accelerator.v:3616" *)
  wire _T_267;
  (* src = "crypto_accelerator.v:4803" *)
  wire _T_2670;
  (* src = "crypto_accelerator.v:4804" *)
  wire _T_2672;
  (* src = "crypto_accelerator.v:4805" *)
  wire _T_2674;
  (* src = "crypto_accelerator.v:4806" *)
  wire _T_2676;
  (* src = "crypto_accelerator.v:4807" *)
  wire _T_2678;
  (* src = "crypto_accelerator.v:4808" *)
  wire _T_2680;
  (* src = "crypto_accelerator.v:4809" *)
  wire _T_2682;
  (* src = "crypto_accelerator.v:4810" *)
  wire _T_2684;
  (* src = "crypto_accelerator.v:4811" *)
  wire _T_2686;
  (* src = "crypto_accelerator.v:4812" *)
  wire _T_2688;
  (* src = "crypto_accelerator.v:3617" *)
  wire _T_269;
  (* src = "crypto_accelerator.v:4813" *)
  wire _T_2690;
  (* src = "crypto_accelerator.v:4814" *)
  wire _T_2692;
  (* src = "crypto_accelerator.v:4815" *)
  wire _T_2694;
  (* src = "crypto_accelerator.v:4816" *)
  wire _T_2696;
  (* src = "crypto_accelerator.v:4817" *)
  wire _T_2698;
  (* src = "crypto_accelerator.v:4818" *)
  wire _T_2700;
  (* src = "crypto_accelerator.v:4819" *)
  wire _T_2702;
  (* src = "crypto_accelerator.v:4820" *)
  wire _T_2704;
  (* src = "crypto_accelerator.v:4821" *)
  wire _T_2706;
  (* src = "crypto_accelerator.v:4822" *)
  wire _T_2708;
  (* src = "crypto_accelerator.v:3618" *)
  wire _T_271;
  (* src = "crypto_accelerator.v:4823" *)
  wire _T_2710;
  (* src = "crypto_accelerator.v:4824" *)
  wire _T_2712;
  (* src = "crypto_accelerator.v:4825" *)
  wire _T_2714;
  (* src = "crypto_accelerator.v:4826" *)
  wire _T_2716;
  (* src = "crypto_accelerator.v:4827" *)
  wire _T_2718;
  (* src = "crypto_accelerator.v:4828" *)
  wire _T_2720;
  (* src = "crypto_accelerator.v:4829" *)
  wire _T_2722;
  (* src = "crypto_accelerator.v:4830" *)
  wire _T_2724;
  (* src = "crypto_accelerator.v:4831" *)
  wire _T_2726;
  (* src = "crypto_accelerator.v:4832" *)
  wire _T_2728;
  (* src = "crypto_accelerator.v:3619" *)
  wire _T_273;
  (* src = "crypto_accelerator.v:4833" *)
  wire _T_2730;
  (* src = "crypto_accelerator.v:4834" *)
  wire _T_2732;
  (* src = "crypto_accelerator.v:4835" *)
  wire _T_2734;
  (* src = "crypto_accelerator.v:4836" *)
  wire _T_2736;
  (* src = "crypto_accelerator.v:4837" *)
  wire _T_2738;
  (* src = "crypto_accelerator.v:4838" *)
  wire _T_2740;
  (* src = "crypto_accelerator.v:4839" *)
  wire _T_2742;
  (* src = "crypto_accelerator.v:4840" *)
  wire _T_2744;
  (* src = "crypto_accelerator.v:4841" *)
  wire _T_2746;
  (* src = "crypto_accelerator.v:4842" *)
  wire _T_2748;
  (* src = "crypto_accelerator.v:3620" *)
  wire _T_275;
  (* src = "crypto_accelerator.v:4843" *)
  wire _T_2750;
  (* src = "crypto_accelerator.v:4844" *)
  wire _T_2752;
  (* src = "crypto_accelerator.v:4845" *)
  wire _T_2754;
  (* src = "crypto_accelerator.v:4846" *)
  wire _T_2756;
  (* src = "crypto_accelerator.v:4847" *)
  wire _T_2758;
  (* src = "crypto_accelerator.v:4848" *)
  wire _T_2760;
  (* src = "crypto_accelerator.v:4849" *)
  wire _T_2762;
  (* src = "crypto_accelerator.v:4850" *)
  wire _T_2764;
  (* src = "crypto_accelerator.v:4851" *)
  wire _T_2766;
  (* src = "crypto_accelerator.v:4852" *)
  wire _T_2768;
  (* src = "crypto_accelerator.v:3621" *)
  wire _T_277;
  (* src = "crypto_accelerator.v:4853" *)
  wire _T_2770;
  (* src = "crypto_accelerator.v:4854" *)
  wire _T_2772;
  (* src = "crypto_accelerator.v:4855" *)
  wire _T_2774;
  (* src = "crypto_accelerator.v:4856" *)
  wire _T_2776;
  (* src = "crypto_accelerator.v:4857" *)
  wire _T_2778;
  (* src = "crypto_accelerator.v:4858" *)
  wire _T_2780;
  (* src = "crypto_accelerator.v:4859" *)
  wire _T_2782;
  (* src = "crypto_accelerator.v:4860" *)
  wire _T_2784;
  (* src = "crypto_accelerator.v:4861" *)
  wire _T_2786;
  (* src = "crypto_accelerator.v:4862" *)
  wire _T_2788;
  (* src = "crypto_accelerator.v:3622" *)
  wire _T_279;
  (* src = "crypto_accelerator.v:4863" *)
  wire _T_2790;
  (* src = "crypto_accelerator.v:4864" *)
  wire _T_2792;
  (* src = "crypto_accelerator.v:4865" *)
  wire _T_2794;
  (* src = "crypto_accelerator.v:4866" *)
  wire _T_2796;
  (* src = "crypto_accelerator.v:4867" *)
  wire _T_2798;
  (* src = "crypto_accelerator.v:4868" *)
  wire _T_2800;
  (* src = "crypto_accelerator.v:4869" *)
  wire _T_2801;
  (* src = "crypto_accelerator.v:4870" *)
  wire _T_2802;
  (* src = "crypto_accelerator.v:4871" *)
  wire _T_2803;
  (* src = "crypto_accelerator.v:4872" *)
  wire _T_2804;
  (* src = "crypto_accelerator.v:4873" *)
  wire _T_2805;
  (* src = "crypto_accelerator.v:4874" *)
  wire _T_2806;
  (* src = "crypto_accelerator.v:4875" *)
  wire _T_2807;
  (* src = "crypto_accelerator.v:4876" *)
  wire _T_2808;
  (* src = "crypto_accelerator.v:3623" *)
  wire _T_281;
  (* src = "crypto_accelerator.v:3624" *)
  wire _T_283;
  (* src = "crypto_accelerator.v:4878" *)
  wire _T_2833;
  (* src = "crypto_accelerator.v:4879" *)
  wire _T_2835;
  (* src = "crypto_accelerator.v:4880" *)
  wire _T_2836;
  (* src = "crypto_accelerator.v:4881" *)
  wire _T_2838;
  (* src = "crypto_accelerator.v:4882" *)
  wire _T_2839;
  (* src = "crypto_accelerator.v:4883" *)
  wire _T_2841;
  (* src = "crypto_accelerator.v:4884" *)
  wire _T_2843;
  (* src = "crypto_accelerator.v:4885" *)
  wire _T_2844;
  (* src = "crypto_accelerator.v:4886" *)
  wire _T_2846;
  (* src = "crypto_accelerator.v:4887" *)
  wire _T_2848;
  (* src = "crypto_accelerator.v:4888" *)
  wire _T_2849;
  (* src = "crypto_accelerator.v:3625" *)
  wire _T_285;
  (* src = "crypto_accelerator.v:4889" *)
  wire _T_2851;
  (* src = "crypto_accelerator.v:4890" *)
  wire _T_2853;
  (* src = "crypto_accelerator.v:4891" *)
  wire _T_2854;
  (* src = "crypto_accelerator.v:4892" *)
  wire _T_2856;
  (* src = "crypto_accelerator.v:4893" *)
  wire _T_2858;
  (* src = "crypto_accelerator.v:4894" *)
  wire _T_2860;
  (* src = "crypto_accelerator.v:4895" *)
  wire _T_2862;
  (* src = "crypto_accelerator.v:4896" *)
  wire _T_2863;
  (* src = "crypto_accelerator.v:4897" *)
  wire _T_2865;
  (* src = "crypto_accelerator.v:4898" *)
  wire _T_2867;
  (* src = "crypto_accelerator.v:4899" *)
  wire _T_2868;
  (* src = "crypto_accelerator.v:3626" *)
  wire _T_287;
  (* src = "crypto_accelerator.v:4900" *)
  wire _T_2870;
  (* src = "crypto_accelerator.v:4901" *)
  wire _T_2872;
  (* src = "crypto_accelerator.v:4902" *)
  wire _T_2874;
  (* src = "crypto_accelerator.v:4903" *)
  wire _T_2875;
  (* src = "crypto_accelerator.v:4904" *)
  wire _T_2877;
  (* src = "crypto_accelerator.v:4905" *)
  wire _T_2878;
  (* src = "crypto_accelerator.v:3627" *)
  wire _T_288;
  (* src = "crypto_accelerator.v:4906" *)
  wire _T_2880;
  (* src = "crypto_accelerator.v:4907" *)
  wire _T_2881;
  (* src = "crypto_accelerator.v:4908" *)
  wire _T_2883;
  (* src = "crypto_accelerator.v:4909" *)
  wire _T_2885;
  (* src = "crypto_accelerator.v:4910" *)
  wire _T_2887;
  (* src = "crypto_accelerator.v:4911" *)
  wire _T_2889;
  (* src = "crypto_accelerator.v:3628" *)
  wire _T_289;
  (* src = "crypto_accelerator.v:4912" *)
  wire _T_2891;
  (* src = "crypto_accelerator.v:4913" *)
  wire _T_2893;
  (* src = "crypto_accelerator.v:4914" *)
  wire _T_2895;
  (* src = "crypto_accelerator.v:4915" *)
  wire _T_2897;
  (* src = "crypto_accelerator.v:4916" *)
  wire _T_2899;
  (* src = "crypto_accelerator.v:3629" *)
  wire _T_290;
  (* src = "crypto_accelerator.v:4917" *)
  wire _T_2901;
  (* src = "crypto_accelerator.v:4918" *)
  wire _T_2903;
  (* src = "crypto_accelerator.v:4919" *)
  wire _T_2905;
  (* src = "crypto_accelerator.v:4920" *)
  wire _T_2907;
  (* src = "crypto_accelerator.v:4921" *)
  wire _T_2909;
  (* src = "crypto_accelerator.v:3630" *)
  wire _T_291;
  (* src = "crypto_accelerator.v:4922" *)
  wire _T_2911;
  (* src = "crypto_accelerator.v:4923" *)
  wire _T_2913;
  (* src = "crypto_accelerator.v:4924" *)
  wire _T_2915;
  (* src = "crypto_accelerator.v:4925" *)
  wire _T_2917;
  (* src = "crypto_accelerator.v:4926" *)
  wire _T_2919;
  (* src = "crypto_accelerator.v:3631" *)
  wire _T_292;
  (* src = "crypto_accelerator.v:4927" *)
  wire _T_2921;
  (* src = "crypto_accelerator.v:4928" *)
  wire _T_2923;
  (* src = "crypto_accelerator.v:4929" *)
  wire _T_2925;
  (* src = "crypto_accelerator.v:4930" *)
  wire _T_2927;
  (* src = "crypto_accelerator.v:4931" *)
  wire _T_2929;
  (* src = "crypto_accelerator.v:3632" *)
  wire _T_293;
  (* src = "crypto_accelerator.v:4932" *)
  wire _T_2931;
  (* src = "crypto_accelerator.v:4933" *)
  wire _T_2933;
  (* src = "crypto_accelerator.v:4934" *)
  wire _T_2935;
  (* src = "crypto_accelerator.v:4935" *)
  wire _T_2937;
  (* src = "crypto_accelerator.v:4936" *)
  wire _T_2939;
  (* src = "crypto_accelerator.v:3633" *)
  wire _T_294;
  (* src = "crypto_accelerator.v:4937" *)
  wire _T_2941;
  (* src = "crypto_accelerator.v:4938" *)
  wire _T_2943;
  (* src = "crypto_accelerator.v:4939" *)
  wire _T_2945;
  (* src = "crypto_accelerator.v:4940" *)
  wire _T_2947;
  (* src = "crypto_accelerator.v:4941" *)
  wire _T_2949;
  (* src = "crypto_accelerator.v:3634" *)
  wire _T_295;
  (* src = "crypto_accelerator.v:4942" *)
  wire _T_2951;
  (* src = "crypto_accelerator.v:4943" *)
  wire _T_2953;
  (* src = "crypto_accelerator.v:4944" *)
  wire _T_2955;
  (* src = "crypto_accelerator.v:4945" *)
  wire _T_2957;
  (* src = "crypto_accelerator.v:4946" *)
  wire _T_2959;
  (* src = "crypto_accelerator.v:4947" *)
  wire _T_2961;
  (* src = "crypto_accelerator.v:4948" *)
  wire _T_2963;
  (* src = "crypto_accelerator.v:4949" *)
  wire _T_2965;
  (* src = "crypto_accelerator.v:4950" *)
  wire _T_2967;
  (* src = "crypto_accelerator.v:4951" *)
  wire _T_2969;
  (* src = "crypto_accelerator.v:4952" *)
  wire _T_2971;
  (* src = "crypto_accelerator.v:4953" *)
  wire _T_2973;
  (* src = "crypto_accelerator.v:4954" *)
  wire _T_2975;
  (* src = "crypto_accelerator.v:4955" *)
  wire _T_2977;
  (* src = "crypto_accelerator.v:4956" *)
  wire _T_2979;
  (* src = "crypto_accelerator.v:4957" *)
  wire _T_2981;
  (* src = "crypto_accelerator.v:4958" *)
  wire _T_2983;
  (* src = "crypto_accelerator.v:4959" *)
  wire _T_2985;
  (* src = "crypto_accelerator.v:4960" *)
  wire _T_2987;
  (* src = "crypto_accelerator.v:4961" *)
  wire _T_2989;
  (* src = "crypto_accelerator.v:4962" *)
  wire _T_2991;
  (* src = "crypto_accelerator.v:4963" *)
  wire _T_2993;
  (* src = "crypto_accelerator.v:4964" *)
  wire _T_2995;
  (* src = "crypto_accelerator.v:4965" *)
  wire _T_2997;
  (* src = "crypto_accelerator.v:4966" *)
  wire _T_2999;
  (* src = "crypto_accelerator.v:4967" *)
  wire _T_3001;
  (* src = "crypto_accelerator.v:4968" *)
  wire _T_3003;
  (* src = "crypto_accelerator.v:4969" *)
  wire _T_3005;
  (* src = "crypto_accelerator.v:4970" *)
  wire _T_3007;
  (* src = "crypto_accelerator.v:4971" *)
  wire _T_3009;
  (* src = "crypto_accelerator.v:4972" *)
  wire _T_3011;
  (* src = "crypto_accelerator.v:4973" *)
  wire _T_3013;
  (* src = "crypto_accelerator.v:4974" *)
  wire _T_3015;
  (* src = "crypto_accelerator.v:4975" *)
  wire _T_3017;
  (* src = "crypto_accelerator.v:4976" *)
  wire _T_3019;
  (* src = "crypto_accelerator.v:4977" *)
  wire _T_3021;
  (* src = "crypto_accelerator.v:4978" *)
  wire _T_3023;
  (* src = "crypto_accelerator.v:4979" *)
  wire _T_3025;
  (* src = "crypto_accelerator.v:4980" *)
  wire _T_3027;
  (* src = "crypto_accelerator.v:4981" *)
  wire _T_3029;
  (* src = "crypto_accelerator.v:4982" *)
  wire _T_3031;
  (* src = "crypto_accelerator.v:4983" *)
  wire _T_3033;
  (* src = "crypto_accelerator.v:4984" *)
  wire _T_3035;
  (* src = "crypto_accelerator.v:4985" *)
  wire _T_3037;
  (* src = "crypto_accelerator.v:4986" *)
  wire _T_3039;
  (* src = "crypto_accelerator.v:4987" *)
  wire _T_3041;
  (* src = "crypto_accelerator.v:4988" *)
  wire _T_3043;
  (* src = "crypto_accelerator.v:4989" *)
  wire _T_3045;
  (* src = "crypto_accelerator.v:4990" *)
  wire _T_3047;
  (* src = "crypto_accelerator.v:4991" *)
  wire _T_3049;
  (* src = "crypto_accelerator.v:4992" *)
  wire _T_3051;
  (* src = "crypto_accelerator.v:4993" *)
  wire _T_3053;
  (* src = "crypto_accelerator.v:4994" *)
  wire _T_3055;
  (* src = "crypto_accelerator.v:4995" *)
  wire _T_3057;
  (* src = "crypto_accelerator.v:4996" *)
  wire _T_3059;
  (* src = "crypto_accelerator.v:4997" *)
  wire _T_3061;
  (* src = "crypto_accelerator.v:4998" *)
  wire _T_3063;
  (* src = "crypto_accelerator.v:4999" *)
  wire _T_3065;
  (* src = "crypto_accelerator.v:5000" *)
  wire _T_3067;
  (* src = "crypto_accelerator.v:5001" *)
  wire _T_3069;
  (* src = "crypto_accelerator.v:5002" *)
  wire _T_3071;
  (* src = "crypto_accelerator.v:5003" *)
  wire _T_3073;
  (* src = "crypto_accelerator.v:5004" *)
  wire _T_3075;
  (* src = "crypto_accelerator.v:5005" *)
  wire _T_3077;
  (* src = "crypto_accelerator.v:5006" *)
  wire _T_3079;
  (* src = "crypto_accelerator.v:5007" *)
  wire _T_3080;
  (* src = "crypto_accelerator.v:5008" *)
  wire _T_3081;
  (* src = "crypto_accelerator.v:5009" *)
  wire _T_3082;
  (* src = "crypto_accelerator.v:5010" *)
  wire _T_3083;
  (* src = "crypto_accelerator.v:5011" *)
  wire _T_3084;
  (* src = "crypto_accelerator.v:5012" *)
  wire _T_3085;
  (* src = "crypto_accelerator.v:5013" *)
  wire _T_3086;
  (* src = "crypto_accelerator.v:5014" *)
  wire _T_3087;
  (* src = "crypto_accelerator.v:5016" *)
  wire _T_3112;
  (* src = "crypto_accelerator.v:5017" *)
  wire _T_3114;
  (* src = "crypto_accelerator.v:5018" *)
  wire _T_3115;
  (* src = "crypto_accelerator.v:5019" *)
  wire _T_3117;
  (* src = "crypto_accelerator.v:5020" *)
  wire _T_3118;
  (* src = "crypto_accelerator.v:5021" *)
  wire _T_3120;
  (* src = "crypto_accelerator.v:5022" *)
  wire _T_3122;
  (* src = "crypto_accelerator.v:5023" *)
  wire _T_3123;
  (* src = "crypto_accelerator.v:5024" *)
  wire _T_3125;
  (* src = "crypto_accelerator.v:5025" *)
  wire _T_3127;
  (* src = "crypto_accelerator.v:5026" *)
  wire _T_3128;
  (* src = "crypto_accelerator.v:5027" *)
  wire _T_3130;
  (* src = "crypto_accelerator.v:5028" *)
  wire _T_3132;
  (* src = "crypto_accelerator.v:5029" *)
  wire _T_3133;
  (* src = "crypto_accelerator.v:5030" *)
  wire _T_3135;
  (* src = "crypto_accelerator.v:5031" *)
  wire _T_3137;
  (* src = "crypto_accelerator.v:5032" *)
  wire _T_3139;
  (* src = "crypto_accelerator.v:5033" *)
  wire _T_3141;
  (* src = "crypto_accelerator.v:5034" *)
  wire _T_3142;
  (* src = "crypto_accelerator.v:5035" *)
  wire _T_3144;
  (* src = "crypto_accelerator.v:5036" *)
  wire _T_3146;
  (* src = "crypto_accelerator.v:5037" *)
  wire _T_3147;
  (* src = "crypto_accelerator.v:5038" *)
  wire _T_3149;
  (* src = "crypto_accelerator.v:5039" *)
  wire _T_3151;
  (* src = "crypto_accelerator.v:5040" *)
  wire _T_3153;
  (* src = "crypto_accelerator.v:5041" *)
  wire _T_3154;
  (* src = "crypto_accelerator.v:5042" *)
  wire _T_3156;
  (* src = "crypto_accelerator.v:5043" *)
  wire _T_3157;
  (* src = "crypto_accelerator.v:5044" *)
  wire _T_3159;
  (* src = "crypto_accelerator.v:5045" *)
  wire _T_3160;
  (* src = "crypto_accelerator.v:5046" *)
  wire _T_3162;
  (* src = "crypto_accelerator.v:5047" *)
  wire _T_3164;
  (* src = "crypto_accelerator.v:5048" *)
  wire _T_3166;
  (* src = "crypto_accelerator.v:5049" *)
  wire _T_3168;
  (* src = "crypto_accelerator.v:5050" *)
  wire _T_3170;
  (* src = "crypto_accelerator.v:5051" *)
  wire _T_3172;
  (* src = "crypto_accelerator.v:5052" *)
  wire _T_3174;
  (* src = "crypto_accelerator.v:5053" *)
  wire _T_3176;
  (* src = "crypto_accelerator.v:5054" *)
  wire _T_3178;
  (* src = "crypto_accelerator.v:5055" *)
  wire _T_3180;
  (* src = "crypto_accelerator.v:5056" *)
  wire _T_3182;
  (* src = "crypto_accelerator.v:5057" *)
  wire _T_3184;
  (* src = "crypto_accelerator.v:5058" *)
  wire _T_3186;
  (* src = "crypto_accelerator.v:5059" *)
  wire _T_3188;
  (* src = "crypto_accelerator.v:5060" *)
  wire _T_3190;
  (* src = "crypto_accelerator.v:5061" *)
  wire _T_3192;
  (* src = "crypto_accelerator.v:5062" *)
  wire _T_3194;
  (* src = "crypto_accelerator.v:5063" *)
  wire _T_3196;
  (* src = "crypto_accelerator.v:5064" *)
  wire _T_3198;
  (* src = "crypto_accelerator.v:3636" *)
  wire _T_320;
  (* src = "crypto_accelerator.v:5065" *)
  wire _T_3200;
  (* src = "crypto_accelerator.v:5066" *)
  wire _T_3202;
  (* src = "crypto_accelerator.v:5067" *)
  wire _T_3204;
  (* src = "crypto_accelerator.v:5068" *)
  wire _T_3206;
  (* src = "crypto_accelerator.v:5069" *)
  wire _T_3208;
  (* src = "crypto_accelerator.v:5070" *)
  wire _T_3210;
  (* src = "crypto_accelerator.v:5071" *)
  wire _T_3212;
  (* src = "crypto_accelerator.v:5072" *)
  wire _T_3214;
  (* src = "crypto_accelerator.v:5073" *)
  wire _T_3216;
  (* src = "crypto_accelerator.v:5074" *)
  wire _T_3218;
  (* src = "crypto_accelerator.v:3637" *)
  wire _T_322;
  (* src = "crypto_accelerator.v:5075" *)
  wire _T_3220;
  (* src = "crypto_accelerator.v:5076" *)
  wire _T_3222;
  (* src = "crypto_accelerator.v:5077" *)
  wire _T_3224;
  (* src = "crypto_accelerator.v:5078" *)
  wire _T_3226;
  (* src = "crypto_accelerator.v:5079" *)
  wire _T_3228;
  (* src = "crypto_accelerator.v:3638" *)
  wire _T_323;
  (* src = "crypto_accelerator.v:5080" *)
  wire _T_3230;
  (* src = "crypto_accelerator.v:5081" *)
  wire _T_3232;
  (* src = "crypto_accelerator.v:5082" *)
  wire _T_3234;
  (* src = "crypto_accelerator.v:5083" *)
  wire _T_3236;
  (* src = "crypto_accelerator.v:5084" *)
  wire _T_3238;
  (* src = "crypto_accelerator.v:5085" *)
  wire _T_3240;
  (* src = "crypto_accelerator.v:5086" *)
  wire _T_3242;
  (* src = "crypto_accelerator.v:5087" *)
  wire _T_3244;
  (* src = "crypto_accelerator.v:5088" *)
  wire _T_3246;
  (* src = "crypto_accelerator.v:5089" *)
  wire _T_3248;
  (* src = "crypto_accelerator.v:3639" *)
  wire _T_325;
  (* src = "crypto_accelerator.v:5090" *)
  wire _T_3250;
  (* src = "crypto_accelerator.v:5091" *)
  wire _T_3252;
  (* src = "crypto_accelerator.v:5092" *)
  wire _T_3254;
  (* src = "crypto_accelerator.v:5093" *)
  wire _T_3256;
  (* src = "crypto_accelerator.v:5094" *)
  wire _T_3258;
  (* src = "crypto_accelerator.v:3640" *)
  wire _T_326;
  (* src = "crypto_accelerator.v:5095" *)
  wire _T_3260;
  (* src = "crypto_accelerator.v:5096" *)
  wire _T_3262;
  (* src = "crypto_accelerator.v:5097" *)
  wire _T_3264;
  (* src = "crypto_accelerator.v:5098" *)
  wire _T_3266;
  (* src = "crypto_accelerator.v:5099" *)
  wire _T_3268;
  (* src = "crypto_accelerator.v:5100" *)
  wire _T_3270;
  (* src = "crypto_accelerator.v:5101" *)
  wire _T_3272;
  (* src = "crypto_accelerator.v:5102" *)
  wire _T_3274;
  (* src = "crypto_accelerator.v:5103" *)
  wire _T_3276;
  (* src = "crypto_accelerator.v:5104" *)
  wire _T_3278;
  (* src = "crypto_accelerator.v:3641" *)
  wire _T_328;
  (* src = "crypto_accelerator.v:5105" *)
  wire _T_3280;
  (* src = "crypto_accelerator.v:5106" *)
  wire _T_3282;
  (* src = "crypto_accelerator.v:5107" *)
  wire _T_3284;
  (* src = "crypto_accelerator.v:5108" *)
  wire _T_3286;
  (* src = "crypto_accelerator.v:5109" *)
  wire _T_3288;
  (* src = "crypto_accelerator.v:5110" *)
  wire _T_3290;
  (* src = "crypto_accelerator.v:5111" *)
  wire _T_3292;
  (* src = "crypto_accelerator.v:5112" *)
  wire _T_3294;
  (* src = "crypto_accelerator.v:5113" *)
  wire _T_3296;
  (* src = "crypto_accelerator.v:5114" *)
  wire _T_3298;
  (* src = "crypto_accelerator.v:3642" *)
  wire _T_330;
  (* src = "crypto_accelerator.v:5115" *)
  wire _T_3300;
  (* src = "crypto_accelerator.v:5116" *)
  wire _T_3302;
  (* src = "crypto_accelerator.v:5117" *)
  wire _T_3304;
  (* src = "crypto_accelerator.v:5118" *)
  wire _T_3306;
  (* src = "crypto_accelerator.v:5119" *)
  wire _T_3308;
  (* src = "crypto_accelerator.v:3643" *)
  wire _T_331;
  (* src = "crypto_accelerator.v:5120" *)
  wire _T_3310;
  (* src = "crypto_accelerator.v:5121" *)
  wire _T_3312;
  (* src = "crypto_accelerator.v:5122" *)
  wire _T_3314;
  (* src = "crypto_accelerator.v:5123" *)
  wire _T_3316;
  (* src = "crypto_accelerator.v:5124" *)
  wire _T_3318;
  (* src = "crypto_accelerator.v:5125" *)
  wire _T_3320;
  (* src = "crypto_accelerator.v:5126" *)
  wire _T_3322;
  (* src = "crypto_accelerator.v:5127" *)
  wire _T_3324;
  (* src = "crypto_accelerator.v:5128" *)
  wire _T_3326;
  (* src = "crypto_accelerator.v:5129" *)
  wire _T_3328;
  (* src = "crypto_accelerator.v:3644" *)
  wire _T_333;
  (* src = "crypto_accelerator.v:5130" *)
  wire _T_3330;
  (* src = "crypto_accelerator.v:5131" *)
  wire _T_3332;
  (* src = "crypto_accelerator.v:5132" *)
  wire _T_3334;
  (* src = "crypto_accelerator.v:5133" *)
  wire _T_3336;
  (* src = "crypto_accelerator.v:5134" *)
  wire _T_3338;
  (* src = "crypto_accelerator.v:5135" *)
  wire _T_3340;
  (* src = "crypto_accelerator.v:5136" *)
  wire _T_3342;
  (* src = "crypto_accelerator.v:5137" *)
  wire _T_3344;
  (* src = "crypto_accelerator.v:5138" *)
  wire _T_3346;
  (* src = "crypto_accelerator.v:5139" *)
  wire _T_3348;
  (* src = "crypto_accelerator.v:3645" *)
  wire _T_335;
  (* src = "crypto_accelerator.v:5140" *)
  wire _T_3350;
  (* src = "crypto_accelerator.v:5141" *)
  wire _T_3352;
  (* src = "crypto_accelerator.v:5142" *)
  wire _T_3354;
  (* src = "crypto_accelerator.v:5143" *)
  wire _T_3356;
  (* src = "crypto_accelerator.v:5144" *)
  wire _T_3358;
  (* src = "crypto_accelerator.v:5145" *)
  wire _T_3359;
  (* src = "crypto_accelerator.v:3646" *)
  wire _T_336;
  (* src = "crypto_accelerator.v:5146" *)
  wire _T_3360;
  (* src = "crypto_accelerator.v:5147" *)
  wire _T_3361;
  (* src = "crypto_accelerator.v:5148" *)
  wire _T_3362;
  (* src = "crypto_accelerator.v:5149" *)
  wire _T_3363;
  (* src = "crypto_accelerator.v:5150" *)
  wire _T_3364;
  (* src = "crypto_accelerator.v:5151" *)
  wire _T_3365;
  (* src = "crypto_accelerator.v:5152" *)
  wire _T_3366;
  (* src = "crypto_accelerator.v:3647" *)
  wire _T_338;
  (* src = "crypto_accelerator.v:5154" *)
  wire _T_3392;
  (* src = "crypto_accelerator.v:5155" *)
  wire _T_3394;
  (* src = "crypto_accelerator.v:5156" *)
  wire _T_3395;
  (* src = "crypto_accelerator.v:5157" *)
  wire _T_3397;
  (* src = "crypto_accelerator.v:5158" *)
  wire _T_3398;
  (* src = "crypto_accelerator.v:3648" *)
  wire _T_340;
  (* src = "crypto_accelerator.v:5159" *)
  wire _T_3400;
  (* src = "crypto_accelerator.v:5160" *)
  wire _T_3402;
  (* src = "crypto_accelerator.v:5161" *)
  wire _T_3403;
  (* src = "crypto_accelerator.v:5162" *)
  wire _T_3405;
  (* src = "crypto_accelerator.v:5163" *)
  wire _T_3407;
  (* src = "crypto_accelerator.v:5164" *)
  wire _T_3408;
  (* src = "crypto_accelerator.v:3649" *)
  wire _T_341;
  (* src = "crypto_accelerator.v:5165" *)
  wire _T_3410;
  (* src = "crypto_accelerator.v:5166" *)
  wire _T_3412;
  (* src = "crypto_accelerator.v:5167" *)
  wire _T_3413;
  (* src = "crypto_accelerator.v:5168" *)
  wire _T_3415;
  (* src = "crypto_accelerator.v:5169" *)
  wire _T_3417;
  (* src = "crypto_accelerator.v:5170" *)
  wire _T_3419;
  (* src = "crypto_accelerator.v:5171" *)
  wire _T_3421;
  (* src = "crypto_accelerator.v:5172" *)
  wire _T_3422;
  (* src = "crypto_accelerator.v:5173" *)
  wire _T_3424;
  (* src = "crypto_accelerator.v:5174" *)
  wire _T_3426;
  (* src = "crypto_accelerator.v:5175" *)
  wire _T_3427;
  (* src = "crypto_accelerator.v:5176" *)
  wire _T_3429;
  (* src = "crypto_accelerator.v:3650" *)
  wire _T_343;
  (* src = "crypto_accelerator.v:5177" *)
  wire _T_3431;
  (* src = "crypto_accelerator.v:5178" *)
  wire _T_3433;
  (* src = "crypto_accelerator.v:5179" *)
  wire _T_3434;
  (* src = "crypto_accelerator.v:5180" *)
  wire _T_3436;
  (* src = "crypto_accelerator.v:5181" *)
  wire _T_3437;
  (* src = "crypto_accelerator.v:5182" *)
  wire _T_3439;
  (* src = "crypto_accelerator.v:5183" *)
  wire _T_3440;
  (* src = "crypto_accelerator.v:5184" *)
  wire _T_3442;
  (* src = "crypto_accelerator.v:5185" *)
  wire _T_3444;
  (* src = "crypto_accelerator.v:5186" *)
  wire _T_3446;
  (* src = "crypto_accelerator.v:5187" *)
  wire _T_3448;
  (* src = "crypto_accelerator.v:3651" *)
  wire _T_345;
  (* src = "crypto_accelerator.v:5188" *)
  wire _T_3450;
  (* src = "crypto_accelerator.v:5189" *)
  wire _T_3452;
  (* src = "crypto_accelerator.v:5190" *)
  wire _T_3454;
  (* src = "crypto_accelerator.v:5191" *)
  wire _T_3456;
  (* src = "crypto_accelerator.v:5192" *)
  wire _T_3458;
  (* src = "crypto_accelerator.v:5193" *)
  wire _T_3460;
  (* src = "crypto_accelerator.v:5194" *)
  wire _T_3462;
  (* src = "crypto_accelerator.v:5195" *)
  wire _T_3464;
  (* src = "crypto_accelerator.v:5196" *)
  wire _T_3466;
  (* src = "crypto_accelerator.v:5197" *)
  wire _T_3468;
  (* src = "crypto_accelerator.v:3652" *)
  wire _T_347;
  (* src = "crypto_accelerator.v:5198" *)
  wire _T_3470;
  (* src = "crypto_accelerator.v:5199" *)
  wire _T_3472;
  (* src = "crypto_accelerator.v:5200" *)
  wire _T_3474;
  (* src = "crypto_accelerator.v:5201" *)
  wire _T_3476;
  (* src = "crypto_accelerator.v:5202" *)
  wire _T_3478;
  (* src = "crypto_accelerator.v:5203" *)
  wire _T_3480;
  (* src = "crypto_accelerator.v:5204" *)
  wire _T_3482;
  (* src = "crypto_accelerator.v:5205" *)
  wire _T_3484;
  (* src = "crypto_accelerator.v:5206" *)
  wire _T_3486;
  (* src = "crypto_accelerator.v:5207" *)
  wire _T_3488;
  (* src = "crypto_accelerator.v:3653" *)
  wire _T_349;
  (* src = "crypto_accelerator.v:5208" *)
  wire _T_3490;
  (* src = "crypto_accelerator.v:5209" *)
  wire _T_3492;
  (* src = "crypto_accelerator.v:5210" *)
  wire _T_3494;
  (* src = "crypto_accelerator.v:5211" *)
  wire _T_3496;
  (* src = "crypto_accelerator.v:5212" *)
  wire _T_3498;
  (* src = "crypto_accelerator.v:3654" *)
  wire _T_350;
  (* src = "crypto_accelerator.v:5213" *)
  wire _T_3500;
  (* src = "crypto_accelerator.v:5214" *)
  wire _T_3502;
  (* src = "crypto_accelerator.v:5215" *)
  wire _T_3504;
  (* src = "crypto_accelerator.v:5216" *)
  wire _T_3506;
  (* src = "crypto_accelerator.v:5217" *)
  wire _T_3508;
  (* src = "crypto_accelerator.v:5218" *)
  wire _T_3510;
  (* src = "crypto_accelerator.v:5219" *)
  wire _T_3512;
  (* src = "crypto_accelerator.v:5220" *)
  wire _T_3514;
  (* src = "crypto_accelerator.v:5221" *)
  wire _T_3516;
  (* src = "crypto_accelerator.v:5222" *)
  wire _T_3518;
  (* src = "crypto_accelerator.v:3655" *)
  wire _T_352;
  (* src = "crypto_accelerator.v:5223" *)
  wire _T_3520;
  (* src = "crypto_accelerator.v:5224" *)
  wire _T_3522;
  (* src = "crypto_accelerator.v:5225" *)
  wire _T_3524;
  (* src = "crypto_accelerator.v:5226" *)
  wire _T_3526;
  (* src = "crypto_accelerator.v:5227" *)
  wire _T_3528;
  (* src = "crypto_accelerator.v:5228" *)
  wire _T_3530;
  (* src = "crypto_accelerator.v:5229" *)
  wire _T_3532;
  (* src = "crypto_accelerator.v:5230" *)
  wire _T_3534;
  (* src = "crypto_accelerator.v:5231" *)
  wire _T_3536;
  (* src = "crypto_accelerator.v:5232" *)
  wire _T_3538;
  (* src = "crypto_accelerator.v:3656" *)
  wire _T_354;
  (* src = "crypto_accelerator.v:5233" *)
  wire _T_3540;
  (* src = "crypto_accelerator.v:5234" *)
  wire _T_3542;
  (* src = "crypto_accelerator.v:5235" *)
  wire _T_3544;
  (* src = "crypto_accelerator.v:5236" *)
  wire _T_3546;
  (* src = "crypto_accelerator.v:5237" *)
  wire _T_3548;
  (* src = "crypto_accelerator.v:3657" *)
  wire _T_355;
  (* src = "crypto_accelerator.v:5238" *)
  wire _T_3550;
  (* src = "crypto_accelerator.v:5239" *)
  wire _T_3552;
  (* src = "crypto_accelerator.v:5240" *)
  wire _T_3554;
  (* src = "crypto_accelerator.v:5241" *)
  wire _T_3556;
  (* src = "crypto_accelerator.v:5242" *)
  wire _T_3558;
  (* src = "crypto_accelerator.v:5243" *)
  wire _T_3560;
  (* src = "crypto_accelerator.v:5244" *)
  wire _T_3562;
  (* src = "crypto_accelerator.v:5245" *)
  wire _T_3564;
  (* src = "crypto_accelerator.v:5246" *)
  wire _T_3566;
  (* src = "crypto_accelerator.v:5247" *)
  wire _T_3568;
  (* src = "crypto_accelerator.v:3658" *)
  wire _T_357;
  (* src = "crypto_accelerator.v:5248" *)
  wire _T_3570;
  (* src = "crypto_accelerator.v:5249" *)
  wire _T_3572;
  (* src = "crypto_accelerator.v:5250" *)
  wire _T_3574;
  (* src = "crypto_accelerator.v:5251" *)
  wire _T_3576;
  (* src = "crypto_accelerator.v:5252" *)
  wire _T_3578;
  (* src = "crypto_accelerator.v:5253" *)
  wire _T_3580;
  (* src = "crypto_accelerator.v:5254" *)
  wire _T_3582;
  (* src = "crypto_accelerator.v:5255" *)
  wire _T_3584;
  (* src = "crypto_accelerator.v:5256" *)
  wire _T_3586;
  (* src = "crypto_accelerator.v:5257" *)
  wire _T_3588;
  (* src = "crypto_accelerator.v:3659" *)
  wire _T_359;
  (* src = "crypto_accelerator.v:5258" *)
  wire _T_3590;
  (* src = "crypto_accelerator.v:5259" *)
  wire _T_3592;
  (* src = "crypto_accelerator.v:5260" *)
  wire _T_3594;
  (* src = "crypto_accelerator.v:5261" *)
  wire _T_3596;
  (* src = "crypto_accelerator.v:5262" *)
  wire _T_3598;
  (* src = "crypto_accelerator.v:5263" *)
  wire _T_3600;
  (* src = "crypto_accelerator.v:5264" *)
  wire _T_3602;
  (* src = "crypto_accelerator.v:5265" *)
  wire _T_3604;
  (* src = "crypto_accelerator.v:5266" *)
  wire _T_3606;
  (* src = "crypto_accelerator.v:5267" *)
  wire _T_3608;
  (* src = "crypto_accelerator.v:3660" *)
  wire _T_361;
  (* src = "crypto_accelerator.v:5268" *)
  wire _T_3610;
  (* src = "crypto_accelerator.v:5269" *)
  wire _T_3612;
  (* src = "crypto_accelerator.v:5270" *)
  wire _T_3614;
  (* src = "crypto_accelerator.v:5271" *)
  wire _T_3616;
  (* src = "crypto_accelerator.v:5272" *)
  wire _T_3618;
  (* src = "crypto_accelerator.v:3661" *)
  wire _T_362;
  (* src = "crypto_accelerator.v:5273" *)
  wire _T_3620;
  (* src = "crypto_accelerator.v:5274" *)
  wire _T_3622;
  (* src = "crypto_accelerator.v:5275" *)
  wire _T_3624;
  (* src = "crypto_accelerator.v:5276" *)
  wire _T_3626;
  (* src = "crypto_accelerator.v:5277" *)
  wire _T_3628;
  (* src = "crypto_accelerator.v:5278" *)
  wire _T_3630;
  (* src = "crypto_accelerator.v:5279" *)
  wire _T_3632;
  (* src = "crypto_accelerator.v:5280" *)
  wire _T_3634;
  (* src = "crypto_accelerator.v:5281" *)
  wire _T_3636;
  (* src = "crypto_accelerator.v:5282" *)
  wire _T_3638;
  (* src = "crypto_accelerator.v:5283" *)
  wire _T_3639;
  (* src = "crypto_accelerator.v:3662" *)
  wire _T_364;
  (* src = "crypto_accelerator.v:5284" *)
  wire _T_3640;
  (* src = "crypto_accelerator.v:5285" *)
  wire _T_3641;
  (* src = "crypto_accelerator.v:5286" *)
  wire _T_3642;
  (* src = "crypto_accelerator.v:5287" *)
  wire _T_3643;
  (* src = "crypto_accelerator.v:5288" *)
  wire _T_3644;
  (* src = "crypto_accelerator.v:5289" *)
  wire _T_3645;
  (* src = "crypto_accelerator.v:5290" *)
  wire _T_3646;
  (* src = "crypto_accelerator.v:3663" *)
  wire _T_365;
  (* src = "crypto_accelerator.v:3664" *)
  wire _T_367;
  (* src = "crypto_accelerator.v:5292" *)
  wire _T_3671;
  (* src = "crypto_accelerator.v:5293" *)
  wire _T_3673;
  (* src = "crypto_accelerator.v:5294" *)
  wire _T_3674;
  (* src = "crypto_accelerator.v:5295" *)
  wire _T_3676;
  (* src = "crypto_accelerator.v:5296" *)
  wire _T_3677;
  (* src = "crypto_accelerator.v:5297" *)
  wire _T_3679;
  (* src = "crypto_accelerator.v:3665" *)
  wire _T_368;
  (* src = "crypto_accelerator.v:5298" *)
  wire _T_3681;
  (* src = "crypto_accelerator.v:5299" *)
  wire _T_3682;
  (* src = "crypto_accelerator.v:5300" *)
  wire _T_3684;
  (* src = "crypto_accelerator.v:5301" *)
  wire _T_3686;
  (* src = "crypto_accelerator.v:5302" *)
  wire _T_3687;
  (* src = "crypto_accelerator.v:5303" *)
  wire _T_3689;
  (* src = "crypto_accelerator.v:5304" *)
  wire _T_3691;
  (* src = "crypto_accelerator.v:5305" *)
  wire _T_3692;
  (* src = "crypto_accelerator.v:5306" *)
  wire _T_3694;
  (* src = "crypto_accelerator.v:5307" *)
  wire _T_3696;
  (* src = "crypto_accelerator.v:5308" *)
  wire _T_3698;
  (* src = "crypto_accelerator.v:3666" *)
  wire _T_370;
  (* src = "crypto_accelerator.v:5309" *)
  wire _T_3700;
  (* src = "crypto_accelerator.v:5310" *)
  wire _T_3701;
  (* src = "crypto_accelerator.v:5311" *)
  wire _T_3703;
  (* src = "crypto_accelerator.v:5312" *)
  wire _T_3705;
  (* src = "crypto_accelerator.v:5313" *)
  wire _T_3706;
  (* src = "crypto_accelerator.v:5314" *)
  wire _T_3708;
  (* src = "crypto_accelerator.v:5315" *)
  wire _T_3710;
  (* src = "crypto_accelerator.v:5316" *)
  wire _T_3712;
  (* src = "crypto_accelerator.v:5317" *)
  wire _T_3713;
  (* src = "crypto_accelerator.v:5318" *)
  wire _T_3715;
  (* src = "crypto_accelerator.v:5319" *)
  wire _T_3716;
  (* src = "crypto_accelerator.v:5320" *)
  wire _T_3718;
  (* src = "crypto_accelerator.v:5321" *)
  wire _T_3719;
  (* src = "crypto_accelerator.v:3667" *)
  wire _T_372;
  (* src = "crypto_accelerator.v:5322" *)
  wire _T_3721;
  (* src = "crypto_accelerator.v:5323" *)
  wire _T_3723;
  (* src = "crypto_accelerator.v:5324" *)
  wire _T_3725;
  (* src = "crypto_accelerator.v:5325" *)
  wire _T_3727;
  (* src = "crypto_accelerator.v:5326" *)
  wire _T_3729;
  (* src = "crypto_accelerator.v:5327" *)
  wire _T_3731;
  (* src = "crypto_accelerator.v:5328" *)
  wire _T_3733;
  (* src = "crypto_accelerator.v:5329" *)
  wire _T_3735;
  (* src = "crypto_accelerator.v:5330" *)
  wire _T_3737;
  (* src = "crypto_accelerator.v:5331" *)
  wire _T_3739;
  (* src = "crypto_accelerator.v:3668" *)
  wire _T_374;
  (* src = "crypto_accelerator.v:5332" *)
  wire _T_3741;
  (* src = "crypto_accelerator.v:5333" *)
  wire _T_3743;
  (* src = "crypto_accelerator.v:5334" *)
  wire _T_3745;
  (* src = "crypto_accelerator.v:5335" *)
  wire _T_3747;
  (* src = "crypto_accelerator.v:5336" *)
  wire _T_3749;
  (* src = "crypto_accelerator.v:5337" *)
  wire _T_3751;
  (* src = "crypto_accelerator.v:5338" *)
  wire _T_3753;
  (* src = "crypto_accelerator.v:5339" *)
  wire _T_3755;
  (* src = "crypto_accelerator.v:5340" *)
  wire _T_3757;
  (* src = "crypto_accelerator.v:5341" *)
  wire _T_3759;
  (* src = "crypto_accelerator.v:3669" *)
  wire _T_376;
  (* src = "crypto_accelerator.v:5342" *)
  wire _T_3761;
  (* src = "crypto_accelerator.v:5343" *)
  wire _T_3763;
  (* src = "crypto_accelerator.v:5344" *)
  wire _T_3765;
  (* src = "crypto_accelerator.v:5345" *)
  wire _T_3767;
  (* src = "crypto_accelerator.v:5346" *)
  wire _T_3769;
  (* src = "crypto_accelerator.v:5347" *)
  wire _T_3771;
  (* src = "crypto_accelerator.v:5348" *)
  wire _T_3773;
  (* src = "crypto_accelerator.v:5349" *)
  wire _T_3775;
  (* src = "crypto_accelerator.v:5350" *)
  wire _T_3777;
  (* src = "crypto_accelerator.v:5351" *)
  wire _T_3779;
  (* src = "crypto_accelerator.v:3670" *)
  wire _T_378;
  (* src = "crypto_accelerator.v:5352" *)
  wire _T_3781;
  (* src = "crypto_accelerator.v:5353" *)
  wire _T_3783;
  (* src = "crypto_accelerator.v:5354" *)
  wire _T_3785;
  (* src = "crypto_accelerator.v:5355" *)
  wire _T_3787;
  (* src = "crypto_accelerator.v:5356" *)
  wire _T_3789;
  (* src = "crypto_accelerator.v:5357" *)
  wire _T_3791;
  (* src = "crypto_accelerator.v:5358" *)
  wire _T_3793;
  (* src = "crypto_accelerator.v:5359" *)
  wire _T_3795;
  (* src = "crypto_accelerator.v:5360" *)
  wire _T_3797;
  (* src = "crypto_accelerator.v:5361" *)
  wire _T_3799;
  (* src = "crypto_accelerator.v:3671" *)
  wire _T_380;
  (* src = "crypto_accelerator.v:5362" *)
  wire _T_3801;
  (* src = "crypto_accelerator.v:5363" *)
  wire _T_3803;
  (* src = "crypto_accelerator.v:5364" *)
  wire _T_3805;
  (* src = "crypto_accelerator.v:5365" *)
  wire _T_3807;
  (* src = "crypto_accelerator.v:5366" *)
  wire _T_3809;
  (* src = "crypto_accelerator.v:5367" *)
  wire _T_3811;
  (* src = "crypto_accelerator.v:5368" *)
  wire _T_3813;
  (* src = "crypto_accelerator.v:5369" *)
  wire _T_3815;
  (* src = "crypto_accelerator.v:5370" *)
  wire _T_3817;
  (* src = "crypto_accelerator.v:5371" *)
  wire _T_3819;
  (* src = "crypto_accelerator.v:3672" *)
  wire _T_382;
  (* src = "crypto_accelerator.v:5372" *)
  wire _T_3821;
  (* src = "crypto_accelerator.v:5373" *)
  wire _T_3823;
  (* src = "crypto_accelerator.v:5374" *)
  wire _T_3825;
  (* src = "crypto_accelerator.v:5375" *)
  wire _T_3827;
  (* src = "crypto_accelerator.v:5376" *)
  wire _T_3829;
  (* src = "crypto_accelerator.v:5377" *)
  wire _T_3831;
  (* src = "crypto_accelerator.v:5378" *)
  wire _T_3833;
  (* src = "crypto_accelerator.v:5379" *)
  wire _T_3835;
  (* src = "crypto_accelerator.v:5380" *)
  wire _T_3837;
  (* src = "crypto_accelerator.v:5381" *)
  wire _T_3839;
  (* src = "crypto_accelerator.v:3673" *)
  wire _T_384;
  (* src = "crypto_accelerator.v:5382" *)
  wire _T_3841;
  (* src = "crypto_accelerator.v:5383" *)
  wire _T_3843;
  (* src = "crypto_accelerator.v:5384" *)
  wire _T_3845;
  (* src = "crypto_accelerator.v:5385" *)
  wire _T_3847;
  (* src = "crypto_accelerator.v:5386" *)
  wire _T_3849;
  (* src = "crypto_accelerator.v:5387" *)
  wire _T_3851;
  (* src = "crypto_accelerator.v:5388" *)
  wire _T_3853;
  (* src = "crypto_accelerator.v:5389" *)
  wire _T_3855;
  (* src = "crypto_accelerator.v:5390" *)
  wire _T_3857;
  (* src = "crypto_accelerator.v:5391" *)
  wire _T_3859;
  (* src = "crypto_accelerator.v:3674" *)
  wire _T_386;
  (* src = "crypto_accelerator.v:5392" *)
  wire _T_3861;
  (* src = "crypto_accelerator.v:5393" *)
  wire _T_3863;
  (* src = "crypto_accelerator.v:5394" *)
  wire _T_3865;
  (* src = "crypto_accelerator.v:5395" *)
  wire _T_3867;
  (* src = "crypto_accelerator.v:5396" *)
  wire _T_3869;
  (* src = "crypto_accelerator.v:5397" *)
  wire _T_3871;
  (* src = "crypto_accelerator.v:5398" *)
  wire _T_3873;
  (* src = "crypto_accelerator.v:5399" *)
  wire _T_3875;
  (* src = "crypto_accelerator.v:5400" *)
  wire _T_3877;
  (* src = "crypto_accelerator.v:5401" *)
  wire _T_3879;
  (* src = "crypto_accelerator.v:3675" *)
  wire _T_388;
  (* src = "crypto_accelerator.v:5402" *)
  wire _T_3881;
  (* src = "crypto_accelerator.v:5403" *)
  wire _T_3883;
  (* src = "crypto_accelerator.v:5404" *)
  wire _T_3885;
  (* src = "crypto_accelerator.v:5405" *)
  wire _T_3887;
  (* src = "crypto_accelerator.v:5406" *)
  wire _T_3889;
  (* src = "crypto_accelerator.v:5407" *)
  wire _T_3891;
  (* src = "crypto_accelerator.v:5408" *)
  wire _T_3893;
  (* src = "crypto_accelerator.v:5409" *)
  wire _T_3895;
  (* src = "crypto_accelerator.v:5410" *)
  wire _T_3897;
  (* src = "crypto_accelerator.v:5411" *)
  wire _T_3899;
  (* src = "crypto_accelerator.v:3676" *)
  wire _T_390;
  (* src = "crypto_accelerator.v:5412" *)
  wire _T_3901;
  (* src = "crypto_accelerator.v:5413" *)
  wire _T_3903;
  (* src = "crypto_accelerator.v:5414" *)
  wire _T_3905;
  (* src = "crypto_accelerator.v:5415" *)
  wire _T_3907;
  (* src = "crypto_accelerator.v:5416" *)
  wire _T_3909;
  (* src = "crypto_accelerator.v:5417" *)
  wire _T_3911;
  (* src = "crypto_accelerator.v:5418" *)
  wire _T_3913;
  (* src = "crypto_accelerator.v:5419" *)
  wire _T_3915;
  (* src = "crypto_accelerator.v:5420" *)
  wire _T_3917;
  (* src = "crypto_accelerator.v:5421" *)
  wire _T_3918;
  (* src = "crypto_accelerator.v:5422" *)
  wire _T_3919;
  (* src = "crypto_accelerator.v:3677" *)
  wire _T_392;
  (* src = "crypto_accelerator.v:5423" *)
  wire _T_3920;
  (* src = "crypto_accelerator.v:5424" *)
  wire _T_3921;
  (* src = "crypto_accelerator.v:5425" *)
  wire _T_3922;
  (* src = "crypto_accelerator.v:5426" *)
  wire _T_3923;
  (* src = "crypto_accelerator.v:5427" *)
  wire _T_3924;
  (* src = "crypto_accelerator.v:5428" *)
  wire _T_3925;
  (* src = "crypto_accelerator.v:3678" *)
  wire _T_394;
  (* src = "crypto_accelerator.v:5430" *)
  wire _T_3950;
  (* src = "crypto_accelerator.v:5431" *)
  wire _T_3952;
  (* src = "crypto_accelerator.v:5432" *)
  wire _T_3953;
  (* src = "crypto_accelerator.v:5433" *)
  wire _T_3955;
  (* src = "crypto_accelerator.v:5434" *)
  wire _T_3956;
  (* src = "crypto_accelerator.v:5435" *)
  wire _T_3958;
  (* src = "crypto_accelerator.v:3679" *)
  wire _T_396;
  (* src = "crypto_accelerator.v:5436" *)
  wire _T_3960;
  (* src = "crypto_accelerator.v:5437" *)
  wire _T_3961;
  (* src = "crypto_accelerator.v:5438" *)
  wire _T_3963;
  (* src = "crypto_accelerator.v:5439" *)
  wire _T_3965;
  (* src = "crypto_accelerator.v:5440" *)
  wire _T_3966;
  (* src = "crypto_accelerator.v:5441" *)
  wire _T_3968;
  (* src = "crypto_accelerator.v:5442" *)
  wire _T_3970;
  (* src = "crypto_accelerator.v:5443" *)
  wire _T_3971;
  (* src = "crypto_accelerator.v:5444" *)
  wire _T_3973;
  (* src = "crypto_accelerator.v:5445" *)
  wire _T_3975;
  (* src = "crypto_accelerator.v:5446" *)
  wire _T_3977;
  (* src = "crypto_accelerator.v:5447" *)
  wire _T_3979;
  (* src = "crypto_accelerator.v:3680" *)
  wire _T_398;
  (* src = "crypto_accelerator.v:5448" *)
  wire _T_3980;
  (* src = "crypto_accelerator.v:5449" *)
  wire _T_3982;
  (* src = "crypto_accelerator.v:5450" *)
  wire _T_3984;
  (* src = "crypto_accelerator.v:5451" *)
  wire _T_3985;
  (* src = "crypto_accelerator.v:5452" *)
  wire _T_3987;
  (* src = "crypto_accelerator.v:5453" *)
  wire _T_3989;
  (* src = "crypto_accelerator.v:5454" *)
  wire _T_3991;
  (* src = "crypto_accelerator.v:5455" *)
  wire _T_3992;
  (* src = "crypto_accelerator.v:5456" *)
  wire _T_3994;
  (* src = "crypto_accelerator.v:5457" *)
  wire _T_3995;
  (* src = "crypto_accelerator.v:5458" *)
  wire _T_3997;
  (* src = "crypto_accelerator.v:5459" *)
  wire _T_3998;
  (* src = "crypto_accelerator.v:3681" *)
  wire _T_400;
  (* src = "crypto_accelerator.v:5460" *)
  wire _T_4000;
  (* src = "crypto_accelerator.v:5461" *)
  wire _T_4002;
  (* src = "crypto_accelerator.v:5462" *)
  wire _T_4004;
  (* src = "crypto_accelerator.v:5463" *)
  wire _T_4006;
  (* src = "crypto_accelerator.v:5464" *)
  wire _T_4008;
  (* src = "crypto_accelerator.v:5465" *)
  wire _T_4010;
  (* src = "crypto_accelerator.v:5466" *)
  wire _T_4012;
  (* src = "crypto_accelerator.v:5467" *)
  wire _T_4014;
  (* src = "crypto_accelerator.v:5468" *)
  wire _T_4016;
  (* src = "crypto_accelerator.v:5469" *)
  wire _T_4018;
  (* src = "crypto_accelerator.v:3682" *)
  wire _T_402;
  (* src = "crypto_accelerator.v:5470" *)
  wire _T_4020;
  (* src = "crypto_accelerator.v:5471" *)
  wire _T_4022;
  (* src = "crypto_accelerator.v:5472" *)
  wire _T_4024;
  (* src = "crypto_accelerator.v:5473" *)
  wire _T_4026;
  (* src = "crypto_accelerator.v:5474" *)
  wire _T_4028;
  (* src = "crypto_accelerator.v:5475" *)
  wire _T_4030;
  (* src = "crypto_accelerator.v:5476" *)
  wire _T_4032;
  (* src = "crypto_accelerator.v:5477" *)
  wire _T_4034;
  (* src = "crypto_accelerator.v:5478" *)
  wire _T_4036;
  (* src = "crypto_accelerator.v:5479" *)
  wire _T_4038;
  (* src = "crypto_accelerator.v:3683" *)
  wire _T_404;
  (* src = "crypto_accelerator.v:5480" *)
  wire _T_4040;
  (* src = "crypto_accelerator.v:5481" *)
  wire _T_4042;
  (* src = "crypto_accelerator.v:5482" *)
  wire _T_4044;
  (* src = "crypto_accelerator.v:5483" *)
  wire _T_4046;
  (* src = "crypto_accelerator.v:5484" *)
  wire _T_4048;
  (* src = "crypto_accelerator.v:5485" *)
  wire _T_4050;
  (* src = "crypto_accelerator.v:5486" *)
  wire _T_4052;
  (* src = "crypto_accelerator.v:5487" *)
  wire _T_4054;
  (* src = "crypto_accelerator.v:5488" *)
  wire _T_4056;
  (* src = "crypto_accelerator.v:5489" *)
  wire _T_4058;
  (* src = "crypto_accelerator.v:3684" *)
  wire _T_406;
  (* src = "crypto_accelerator.v:5490" *)
  wire _T_4060;
  (* src = "crypto_accelerator.v:5491" *)
  wire _T_4062;
  (* src = "crypto_accelerator.v:5492" *)
  wire _T_4064;
  (* src = "crypto_accelerator.v:5493" *)
  wire _T_4066;
  (* src = "crypto_accelerator.v:5494" *)
  wire _T_4068;
  (* src = "crypto_accelerator.v:5495" *)
  wire _T_4070;
  (* src = "crypto_accelerator.v:5496" *)
  wire _T_4072;
  (* src = "crypto_accelerator.v:5497" *)
  wire _T_4074;
  (* src = "crypto_accelerator.v:5498" *)
  wire _T_4076;
  (* src = "crypto_accelerator.v:5499" *)
  wire _T_4078;
  (* src = "crypto_accelerator.v:3685" *)
  wire _T_408;
  (* src = "crypto_accelerator.v:5500" *)
  wire _T_4080;
  (* src = "crypto_accelerator.v:5501" *)
  wire _T_4082;
  (* src = "crypto_accelerator.v:5502" *)
  wire _T_4084;
  (* src = "crypto_accelerator.v:5503" *)
  wire _T_4086;
  (* src = "crypto_accelerator.v:5504" *)
  wire _T_4088;
  (* src = "crypto_accelerator.v:5505" *)
  wire _T_4090;
  (* src = "crypto_accelerator.v:5506" *)
  wire _T_4092;
  (* src = "crypto_accelerator.v:5507" *)
  wire _T_4094;
  (* src = "crypto_accelerator.v:5508" *)
  wire _T_4096;
  (* src = "crypto_accelerator.v:5509" *)
  wire _T_4098;
  (* src = "crypto_accelerator.v:3498" *)
  wire _T_41;
  (* src = "crypto_accelerator.v:3686" *)
  wire _T_410;
  (* src = "crypto_accelerator.v:5510" *)
  wire _T_4100;
  (* src = "crypto_accelerator.v:5511" *)
  wire _T_4102;
  (* src = "crypto_accelerator.v:5512" *)
  wire _T_4104;
  (* src = "crypto_accelerator.v:5513" *)
  wire _T_4106;
  (* src = "crypto_accelerator.v:5514" *)
  wire _T_4108;
  (* src = "crypto_accelerator.v:5515" *)
  wire _T_4110;
  (* src = "crypto_accelerator.v:5516" *)
  wire _T_4112;
  (* src = "crypto_accelerator.v:5517" *)
  wire _T_4114;
  (* src = "crypto_accelerator.v:5518" *)
  wire _T_4116;
  (* src = "crypto_accelerator.v:5519" *)
  wire _T_4118;
  (* src = "crypto_accelerator.v:3687" *)
  wire _T_412;
  (* src = "crypto_accelerator.v:5520" *)
  wire _T_4120;
  (* src = "crypto_accelerator.v:5521" *)
  wire _T_4122;
  (* src = "crypto_accelerator.v:5522" *)
  wire _T_4124;
  (* src = "crypto_accelerator.v:5523" *)
  wire _T_4126;
  (* src = "crypto_accelerator.v:5524" *)
  wire _T_4128;
  (* src = "crypto_accelerator.v:5525" *)
  wire _T_4130;
  (* src = "crypto_accelerator.v:5526" *)
  wire _T_4132;
  (* src = "crypto_accelerator.v:5527" *)
  wire _T_4134;
  (* src = "crypto_accelerator.v:5528" *)
  wire _T_4136;
  (* src = "crypto_accelerator.v:5529" *)
  wire _T_4138;
  (* src = "crypto_accelerator.v:3688" *)
  wire _T_414;
  (* src = "crypto_accelerator.v:5530" *)
  wire _T_4140;
  (* src = "crypto_accelerator.v:5531" *)
  wire _T_4142;
  (* src = "crypto_accelerator.v:5532" *)
  wire _T_4144;
  (* src = "crypto_accelerator.v:5533" *)
  wire _T_4146;
  (* src = "crypto_accelerator.v:5534" *)
  wire _T_4148;
  (* src = "crypto_accelerator.v:5535" *)
  wire _T_4150;
  (* src = "crypto_accelerator.v:5536" *)
  wire _T_4152;
  (* src = "crypto_accelerator.v:5537" *)
  wire _T_4154;
  (* src = "crypto_accelerator.v:5538" *)
  wire _T_4156;
  (* src = "crypto_accelerator.v:5539" *)
  wire _T_4158;
  (* src = "crypto_accelerator.v:3689" *)
  wire _T_416;
  (* src = "crypto_accelerator.v:5540" *)
  wire _T_4160;
  (* src = "crypto_accelerator.v:5541" *)
  wire _T_4162;
  (* src = "crypto_accelerator.v:5542" *)
  wire _T_4164;
  (* src = "crypto_accelerator.v:5543" *)
  wire _T_4166;
  (* src = "crypto_accelerator.v:5544" *)
  wire _T_4168;
  (* src = "crypto_accelerator.v:5545" *)
  wire _T_4170;
  (* src = "crypto_accelerator.v:5546" *)
  wire _T_4172;
  (* src = "crypto_accelerator.v:5547" *)
  wire _T_4174;
  (* src = "crypto_accelerator.v:5548" *)
  wire _T_4176;
  (* src = "crypto_accelerator.v:5549" *)
  wire _T_4178;
  (* src = "crypto_accelerator.v:3690" *)
  wire _T_418;
  (* src = "crypto_accelerator.v:5550" *)
  wire _T_4180;
  (* src = "crypto_accelerator.v:5551" *)
  wire _T_4182;
  (* src = "crypto_accelerator.v:5552" *)
  wire _T_4184;
  (* src = "crypto_accelerator.v:5553" *)
  wire _T_4186;
  (* src = "crypto_accelerator.v:5554" *)
  wire _T_4188;
  (* src = "crypto_accelerator.v:5555" *)
  wire _T_4190;
  (* src = "crypto_accelerator.v:5556" *)
  wire _T_4192;
  (* src = "crypto_accelerator.v:5557" *)
  wire _T_4194;
  (* src = "crypto_accelerator.v:5558" *)
  wire _T_4196;
  (* src = "crypto_accelerator.v:5559" *)
  wire _T_4197;
  (* src = "crypto_accelerator.v:5560" *)
  wire _T_4198;
  (* src = "crypto_accelerator.v:5561" *)
  wire _T_4199;
  (* src = "crypto_accelerator.v:3691" *)
  wire _T_420;
  (* src = "crypto_accelerator.v:5562" *)
  wire _T_4200;
  (* src = "crypto_accelerator.v:5563" *)
  wire _T_4201;
  (* src = "crypto_accelerator.v:5564" *)
  wire _T_4202;
  (* src = "crypto_accelerator.v:5565" *)
  wire _T_4203;
  (* src = "crypto_accelerator.v:5566" *)
  wire _T_4204;
  (* src = "crypto_accelerator.v:3692" *)
  wire _T_422;
  (* src = "crypto_accelerator.v:5568" *)
  wire _T_4229;
  (* src = "crypto_accelerator.v:5569" *)
  wire _T_4231;
  (* src = "crypto_accelerator.v:5570" *)
  wire _T_4232;
  (* src = "crypto_accelerator.v:5571" *)
  wire _T_4234;
  (* src = "crypto_accelerator.v:5572" *)
  wire _T_4235;
  (* src = "crypto_accelerator.v:5573" *)
  wire _T_4237;
  (* src = "crypto_accelerator.v:5574" *)
  wire _T_4239;
  (* src = "crypto_accelerator.v:3693" *)
  wire _T_424;
  (* src = "crypto_accelerator.v:5575" *)
  wire _T_4240;
  (* src = "crypto_accelerator.v:5576" *)
  wire _T_4242;
  (* src = "crypto_accelerator.v:5577" *)
  wire _T_4244;
  (* src = "crypto_accelerator.v:5578" *)
  wire _T_4245;
  (* src = "crypto_accelerator.v:5579" *)
  wire _T_4247;
  (* src = "crypto_accelerator.v:5580" *)
  wire _T_4249;
  (* src = "crypto_accelerator.v:5581" *)
  wire _T_4250;
  (* src = "crypto_accelerator.v:5582" *)
  wire _T_4252;
  (* src = "crypto_accelerator.v:5583" *)
  wire _T_4254;
  (* src = "crypto_accelerator.v:5584" *)
  wire _T_4256;
  (* src = "crypto_accelerator.v:5585" *)
  wire _T_4258;
  (* src = "crypto_accelerator.v:5586" *)
  wire _T_4259;
  (* src = "crypto_accelerator.v:3694" *)
  wire _T_426;
  (* src = "crypto_accelerator.v:5587" *)
  wire _T_4261;
  (* src = "crypto_accelerator.v:5588" *)
  wire _T_4263;
  (* src = "crypto_accelerator.v:5589" *)
  wire _T_4264;
  (* src = "crypto_accelerator.v:5590" *)
  wire _T_4266;
  (* src = "crypto_accelerator.v:5591" *)
  wire _T_4268;
  (* src = "crypto_accelerator.v:5592" *)
  wire _T_4270;
  (* src = "crypto_accelerator.v:5593" *)
  wire _T_4271;
  (* src = "crypto_accelerator.v:5594" *)
  wire _T_4273;
  (* src = "crypto_accelerator.v:5595" *)
  wire _T_4274;
  (* src = "crypto_accelerator.v:5596" *)
  wire _T_4276;
  (* src = "crypto_accelerator.v:5597" *)
  wire _T_4277;
  (* src = "crypto_accelerator.v:5598" *)
  wire _T_4279;
  (* src = "crypto_accelerator.v:3695" *)
  wire _T_428;
  (* src = "crypto_accelerator.v:5599" *)
  wire _T_4281;
  (* src = "crypto_accelerator.v:5600" *)
  wire _T_4283;
  (* src = "crypto_accelerator.v:5601" *)
  wire _T_4285;
  (* src = "crypto_accelerator.v:5602" *)
  wire _T_4287;
  (* src = "crypto_accelerator.v:5603" *)
  wire _T_4289;
  (* src = "crypto_accelerator.v:5604" *)
  wire _T_4291;
  (* src = "crypto_accelerator.v:5605" *)
  wire _T_4293;
  (* src = "crypto_accelerator.v:5606" *)
  wire _T_4295;
  (* src = "crypto_accelerator.v:5607" *)
  wire _T_4297;
  (* src = "crypto_accelerator.v:5608" *)
  wire _T_4299;
  (* src = "crypto_accelerator.v:3499" *)
  wire _T_43;
  (* src = "crypto_accelerator.v:3696" *)
  wire _T_430;
  (* src = "crypto_accelerator.v:5609" *)
  wire _T_4301;
  (* src = "crypto_accelerator.v:5610" *)
  wire _T_4303;
  (* src = "crypto_accelerator.v:5611" *)
  wire _T_4305;
  (* src = "crypto_accelerator.v:5612" *)
  wire _T_4307;
  (* src = "crypto_accelerator.v:5613" *)
  wire _T_4309;
  (* src = "crypto_accelerator.v:5614" *)
  wire _T_4311;
  (* src = "crypto_accelerator.v:5615" *)
  wire _T_4313;
  (* src = "crypto_accelerator.v:5616" *)
  wire _T_4315;
  (* src = "crypto_accelerator.v:5617" *)
  wire _T_4317;
  (* src = "crypto_accelerator.v:5618" *)
  wire _T_4319;
  (* src = "crypto_accelerator.v:3697" *)
  wire _T_432;
  (* src = "crypto_accelerator.v:5619" *)
  wire _T_4321;
  (* src = "crypto_accelerator.v:5620" *)
  wire _T_4323;
  (* src = "crypto_accelerator.v:5621" *)
  wire _T_4325;
  (* src = "crypto_accelerator.v:5622" *)
  wire _T_4327;
  (* src = "crypto_accelerator.v:5623" *)
  wire _T_4329;
  (* src = "crypto_accelerator.v:5624" *)
  wire _T_4331;
  (* src = "crypto_accelerator.v:5625" *)
  wire _T_4333;
  (* src = "crypto_accelerator.v:5626" *)
  wire _T_4335;
  (* src = "crypto_accelerator.v:5627" *)
  wire _T_4337;
  (* src = "crypto_accelerator.v:5628" *)
  wire _T_4339;
  (* src = "crypto_accelerator.v:3698" *)
  wire _T_434;
  (* src = "crypto_accelerator.v:5629" *)
  wire _T_4341;
  (* src = "crypto_accelerator.v:5630" *)
  wire _T_4343;
  (* src = "crypto_accelerator.v:5631" *)
  wire _T_4345;
  (* src = "crypto_accelerator.v:5632" *)
  wire _T_4347;
  (* src = "crypto_accelerator.v:5633" *)
  wire _T_4349;
  (* src = "crypto_accelerator.v:5634" *)
  wire _T_4351;
  (* src = "crypto_accelerator.v:5635" *)
  wire _T_4353;
  (* src = "crypto_accelerator.v:5636" *)
  wire _T_4355;
  (* src = "crypto_accelerator.v:5637" *)
  wire _T_4357;
  (* src = "crypto_accelerator.v:5638" *)
  wire _T_4359;
  (* src = "crypto_accelerator.v:3699" *)
  wire _T_436;
  (* src = "crypto_accelerator.v:5639" *)
  wire _T_4361;
  (* src = "crypto_accelerator.v:5640" *)
  wire _T_4363;
  (* src = "crypto_accelerator.v:5641" *)
  wire _T_4365;
  (* src = "crypto_accelerator.v:5642" *)
  wire _T_4367;
  (* src = "crypto_accelerator.v:5643" *)
  wire _T_4369;
  (* src = "crypto_accelerator.v:5644" *)
  wire _T_4371;
  (* src = "crypto_accelerator.v:5645" *)
  wire _T_4373;
  (* src = "crypto_accelerator.v:5646" *)
  wire _T_4375;
  (* src = "crypto_accelerator.v:5647" *)
  wire _T_4377;
  (* src = "crypto_accelerator.v:5648" *)
  wire _T_4379;
  (* src = "crypto_accelerator.v:3700" *)
  wire _T_438;
  (* src = "crypto_accelerator.v:5649" *)
  wire _T_4381;
  (* src = "crypto_accelerator.v:5650" *)
  wire _T_4383;
  (* src = "crypto_accelerator.v:5651" *)
  wire _T_4385;
  (* src = "crypto_accelerator.v:5652" *)
  wire _T_4387;
  (* src = "crypto_accelerator.v:5653" *)
  wire _T_4389;
  (* src = "crypto_accelerator.v:5654" *)
  wire _T_4391;
  (* src = "crypto_accelerator.v:5655" *)
  wire _T_4393;
  (* src = "crypto_accelerator.v:5656" *)
  wire _T_4395;
  (* src = "crypto_accelerator.v:5657" *)
  wire _T_4397;
  (* src = "crypto_accelerator.v:5658" *)
  wire _T_4399;
  (* src = "crypto_accelerator.v:3500" *)
  wire _T_44;
  (* src = "crypto_accelerator.v:3701" *)
  wire _T_440;
  (* src = "crypto_accelerator.v:5659" *)
  wire _T_4401;
  (* src = "crypto_accelerator.v:5660" *)
  wire _T_4403;
  (* src = "crypto_accelerator.v:5661" *)
  wire _T_4405;
  (* src = "crypto_accelerator.v:5662" *)
  wire _T_4407;
  (* src = "crypto_accelerator.v:5663" *)
  wire _T_4409;
  (* src = "crypto_accelerator.v:5664" *)
  wire _T_4411;
  (* src = "crypto_accelerator.v:5665" *)
  wire _T_4413;
  (* src = "crypto_accelerator.v:5666" *)
  wire _T_4415;
  (* src = "crypto_accelerator.v:5667" *)
  wire _T_4417;
  (* src = "crypto_accelerator.v:5668" *)
  wire _T_4419;
  (* src = "crypto_accelerator.v:3702" *)
  wire _T_442;
  (* src = "crypto_accelerator.v:5669" *)
  wire _T_4421;
  (* src = "crypto_accelerator.v:5670" *)
  wire _T_4423;
  (* src = "crypto_accelerator.v:5671" *)
  wire _T_4425;
  (* src = "crypto_accelerator.v:5672" *)
  wire _T_4427;
  (* src = "crypto_accelerator.v:5673" *)
  wire _T_4429;
  (* src = "crypto_accelerator.v:5674" *)
  wire _T_4431;
  (* src = "crypto_accelerator.v:5675" *)
  wire _T_4433;
  (* src = "crypto_accelerator.v:5676" *)
  wire _T_4435;
  (* src = "crypto_accelerator.v:5677" *)
  wire _T_4437;
  (* src = "crypto_accelerator.v:5678" *)
  wire _T_4439;
  (* src = "crypto_accelerator.v:3703" *)
  wire _T_444;
  (* src = "crypto_accelerator.v:5679" *)
  wire _T_4441;
  (* src = "crypto_accelerator.v:5680" *)
  wire _T_4443;
  (* src = "crypto_accelerator.v:5681" *)
  wire _T_4445;
  (* src = "crypto_accelerator.v:5682" *)
  wire _T_4447;
  (* src = "crypto_accelerator.v:5683" *)
  wire _T_4449;
  (* src = "crypto_accelerator.v:5684" *)
  wire _T_4451;
  (* src = "crypto_accelerator.v:5685" *)
  wire _T_4453;
  (* src = "crypto_accelerator.v:5686" *)
  wire _T_4455;
  (* src = "crypto_accelerator.v:5687" *)
  wire _T_4457;
  (* src = "crypto_accelerator.v:5688" *)
  wire _T_4459;
  (* src = "crypto_accelerator.v:3704" *)
  wire _T_446;
  (* src = "crypto_accelerator.v:5689" *)
  wire _T_4461;
  (* src = "crypto_accelerator.v:5690" *)
  wire _T_4463;
  (* src = "crypto_accelerator.v:5691" *)
  wire _T_4465;
  (* src = "crypto_accelerator.v:5692" *)
  wire _T_4467;
  (* src = "crypto_accelerator.v:5693" *)
  wire _T_4469;
  (* src = "crypto_accelerator.v:5694" *)
  wire _T_4471;
  (* src = "crypto_accelerator.v:5695" *)
  wire _T_4473;
  (* src = "crypto_accelerator.v:5696" *)
  wire _T_4475;
  (* src = "crypto_accelerator.v:5697" *)
  wire _T_4476;
  (* src = "crypto_accelerator.v:5698" *)
  wire _T_4477;
  (* src = "crypto_accelerator.v:5699" *)
  wire _T_4478;
  (* src = "crypto_accelerator.v:5700" *)
  wire _T_4479;
  (* src = "crypto_accelerator.v:3705" *)
  wire _T_448;
  (* src = "crypto_accelerator.v:5701" *)
  wire _T_4480;
  (* src = "crypto_accelerator.v:5702" *)
  wire _T_4481;
  (* src = "crypto_accelerator.v:5703" *)
  wire _T_4482;
  (* src = "crypto_accelerator.v:5704" *)
  wire _T_4483;
  (* src = "crypto_accelerator.v:3706" *)
  wire _T_450;
  (* src = "crypto_accelerator.v:3707" *)
  wire _T_452;
  (* src = "crypto_accelerator.v:5947" *)
  wire [7:0] _T_4534;
  (* src = "crypto_accelerator.v:5948" *)
  wire [7:0] _T_4535;
  (* src = "crypto_accelerator.v:5949" *)
  wire _T_4536;
  (* src = "crypto_accelerator.v:5950" *)
  wire [8:0] _T_4537;
  (* src = "crypto_accelerator.v:5951" *)
  wire [8:0] _T_4538;
  (* src = "crypto_accelerator.v:5952" *)
  wire [8:0] _T_4539;
  (* src = "crypto_accelerator.v:3708" *)
  wire _T_454;
  (* src = "crypto_accelerator.v:5953" *)
  wire [8:0] _T_4541;
  (* src = "crypto_accelerator.v:5954" *)
  wire [8:0] _T_4542;
  (* src = "crypto_accelerator.v:5955" *)
  wire _T_4543;
  (* src = "crypto_accelerator.v:5956" *)
  wire [9:0] _T_4544;
  wire [7:0] _T_4545;
  wire [7:0] _T_4546;
  wire [7:0] _T_4548;
  (* src = "crypto_accelerator.v:5960" *)
  wire [7:0] _T_4549;
  (* src = "crypto_accelerator.v:5961" *)
  wire [7:0] _T_4550;
  (* src = "crypto_accelerator.v:5962" *)
  wire _T_4551;
  (* src = "crypto_accelerator.v:5963" *)
  wire [8:0] _T_4552;
  (* src = "crypto_accelerator.v:5964" *)
  wire [8:0] _T_4553;
  (* src = "crypto_accelerator.v:5965" *)
  wire [8:0] _T_4554;
  (* src = "crypto_accelerator.v:5966" *)
  wire [8:0] _T_4556;
  (* src = "crypto_accelerator.v:5967" *)
  wire [8:0] _T_4557;
  (* src = "crypto_accelerator.v:5968" *)
  wire _T_4558;
  (* src = "crypto_accelerator.v:5969" *)
  wire [9:0] _T_4559;
  (* src = "crypto_accelerator.v:3709" *)
  wire _T_456;
  wire [7:0] _T_4560;
  wire [7:0] _T_4561;
  wire [7:0] _T_4563;
  (* src = "crypto_accelerator.v:5974" *)
  wire [9:0] _T_4564;
  (* src = "crypto_accelerator.v:5976" *)
  wire [9:0] _T_4565;
  (* src = "crypto_accelerator.v:5978" *)
  wire [9:0] _T_4566;
  (* src = "crypto_accelerator.v:5980" *)
  wire [9:0] _T_4567;
  (* src = "crypto_accelerator.v:5981" *)
  wire [7:0] _T_4568;
  (* src = "crypto_accelerator.v:5982" *)
  wire [7:0] _T_4569;
  (* src = "crypto_accelerator.v:5983" *)
  wire _T_4570;
  (* src = "crypto_accelerator.v:5984" *)
  wire [8:0] _T_4571;
  (* src = "crypto_accelerator.v:5985" *)
  wire [8:0] _T_4572;
  (* src = "crypto_accelerator.v:5986" *)
  wire [8:0] _T_4573;
  (* src = "crypto_accelerator.v:5987" *)
  wire [8:0] _T_4575;
  (* src = "crypto_accelerator.v:5988" *)
  wire [8:0] _T_4576;
  (* src = "crypto_accelerator.v:5989" *)
  wire _T_4577;
  (* src = "crypto_accelerator.v:5990" *)
  wire [9:0] _T_4578;
  wire [7:0] _T_4579;
  (* src = "crypto_accelerator.v:3710" *)
  wire _T_458;
  wire [7:0] _T_4580;
  (* src = "crypto_accelerator.v:5993" *)
  wire [9:0] _T_4582;
  (* src = "crypto_accelerator.v:5994" *)
  wire [7:0] _T_4583;
  (* src = "crypto_accelerator.v:5995" *)
  wire [7:0] _T_4584;
  (* src = "crypto_accelerator.v:5996" *)
  wire _T_4585;
  (* src = "crypto_accelerator.v:5997" *)
  wire [8:0] _T_4586;
  (* src = "crypto_accelerator.v:5998" *)
  wire [8:0] _T_4587;
  (* src = "crypto_accelerator.v:5999" *)
  wire [8:0] _T_4588;
  (* src = "crypto_accelerator.v:6000" *)
  wire [8:0] _T_4590;
  (* src = "crypto_accelerator.v:6001" *)
  wire [8:0] _T_4591;
  (* src = "crypto_accelerator.v:6002" *)
  wire _T_4592;
  (* src = "crypto_accelerator.v:6003" *)
  wire [9:0] _T_4593;
  wire [7:0] _T_4594;
  (* src = "crypto_accelerator.v:6005" *)
  wire [9:0] _T_4595;
  wire [7:0] _T_4597;
  (* src = "crypto_accelerator.v:6008" *)
  wire [9:0] _T_4598;
  (* src = "crypto_accelerator.v:6010" *)
  wire [9:0] _T_4599;
  (* src = "crypto_accelerator.v:3501" *)
  wire _T_46;
  (* src = "crypto_accelerator.v:3711" *)
  wire _T_460;
  (* src = "crypto_accelerator.v:6012" *)
  wire [9:0] _T_4600;
  (* src = "crypto_accelerator.v:6014" *)
  wire [9:0] _T_4601;
  (* src = "crypto_accelerator.v:6015" *)
  wire [7:0] _T_4602;
  (* src = "crypto_accelerator.v:6016" *)
  wire [7:0] _T_4603;
  (* src = "crypto_accelerator.v:6017" *)
  wire _T_4604;
  (* src = "crypto_accelerator.v:6018" *)
  wire [8:0] _T_4605;
  (* src = "crypto_accelerator.v:6019" *)
  wire [8:0] _T_4606;
  (* src = "crypto_accelerator.v:6020" *)
  wire [8:0] _T_4607;
  (* src = "crypto_accelerator.v:6021" *)
  wire [8:0] _T_4609;
  (* src = "crypto_accelerator.v:6022" *)
  wire [8:0] _T_4610;
  (* src = "crypto_accelerator.v:6023" *)
  wire _T_4611;
  (* src = "crypto_accelerator.v:6024" *)
  wire [9:0] _T_4612;
  wire [7:0] _T_4613;
  wire [7:0] _T_4614;
  (* src = "crypto_accelerator.v:6027" *)
  wire [9:0] _T_4616;
  (* src = "crypto_accelerator.v:6028" *)
  wire [7:0] _T_4617;
  (* src = "crypto_accelerator.v:6029" *)
  wire [7:0] _T_4618;
  (* src = "crypto_accelerator.v:6030" *)
  wire _T_4619;
  (* src = "crypto_accelerator.v:3712" *)
  wire _T_462;
  (* src = "crypto_accelerator.v:6031" *)
  wire [8:0] _T_4620;
  (* src = "crypto_accelerator.v:6032" *)
  wire [8:0] _T_4621;
  (* src = "crypto_accelerator.v:6033" *)
  wire [8:0] _T_4622;
  (* src = "crypto_accelerator.v:6034" *)
  wire [8:0] _T_4624;
  (* src = "crypto_accelerator.v:6035" *)
  wire [8:0] _T_4625;
  (* src = "crypto_accelerator.v:6036" *)
  wire _T_4626;
  (* src = "crypto_accelerator.v:6037" *)
  wire [9:0] _T_4627;
  wire [7:0] _T_4628;
  (* src = "crypto_accelerator.v:6039" *)
  wire [9:0] _T_4629;
  (* src = "crypto_accelerator.v:6040" *)
  wire [9:0] _T_4631;
  (* src = "crypto_accelerator.v:6042" *)
  wire [9:0] _T_4632;
  (* src = "crypto_accelerator.v:6044" *)
  wire [9:0] _T_4633;
  (* src = "crypto_accelerator.v:6046" *)
  wire [9:0] _T_4634;
  (* src = "crypto_accelerator.v:6048" *)
  wire [9:0] _T_4635;
  (* src = "crypto_accelerator.v:6049" *)
  wire [7:0] _T_4636;
  (* src = "crypto_accelerator.v:6050" *)
  wire [7:0] _T_4637;
  (* src = "crypto_accelerator.v:6051" *)
  wire _T_4638;
  (* src = "crypto_accelerator.v:6052" *)
  wire [8:0] _T_4639;
  (* src = "crypto_accelerator.v:3713" *)
  wire _T_464;
  (* src = "crypto_accelerator.v:6053" *)
  wire [8:0] _T_4640;
  (* src = "crypto_accelerator.v:6054" *)
  wire [8:0] _T_4641;
  (* src = "crypto_accelerator.v:6055" *)
  wire [8:0] _T_4643;
  (* src = "crypto_accelerator.v:6056" *)
  wire [8:0] _T_4644;
  (* src = "crypto_accelerator.v:6057" *)
  wire _T_4645;
  (* src = "crypto_accelerator.v:6058" *)
  wire [9:0] _T_4646;
  wire [7:0] _T_4647;
  wire [7:0] _T_4648;
  (* src = "crypto_accelerator.v:6061" *)
  wire [9:0] _T_4650;
  (* src = "crypto_accelerator.v:6062" *)
  wire [7:0] _T_4651;
  (* src = "crypto_accelerator.v:6063" *)
  wire [7:0] _T_4652;
  (* src = "crypto_accelerator.v:6064" *)
  wire _T_4653;
  (* src = "crypto_accelerator.v:6065" *)
  wire [8:0] _T_4654;
  (* src = "crypto_accelerator.v:6066" *)
  wire [8:0] _T_4655;
  (* src = "crypto_accelerator.v:6067" *)
  wire [8:0] _T_4656;
  (* src = "crypto_accelerator.v:6068" *)
  wire [8:0] _T_4658;
  (* src = "crypto_accelerator.v:6069" *)
  wire [8:0] _T_4659;
  (* src = "crypto_accelerator.v:3714" *)
  wire _T_466;
  (* src = "crypto_accelerator.v:6070" *)
  wire _T_4660;
  (* src = "crypto_accelerator.v:6071" *)
  wire [9:0] _T_4661;
  wire [7:0] _T_4662;
  (* src = "crypto_accelerator.v:6073" *)
  wire [9:0] _T_4663;
  wire [7:0] _T_4665;
  (* src = "crypto_accelerator.v:6076" *)
  wire [9:0] _T_4666;
  (* src = "crypto_accelerator.v:6078" *)
  wire [9:0] _T_4667;
  (* src = "crypto_accelerator.v:6080" *)
  wire [9:0] _T_4668;
  (* src = "crypto_accelerator.v:6082" *)
  wire [9:0] _T_4669;
  (* src = "crypto_accelerator.v:3715" *)
  wire _T_468;
  (* src = "crypto_accelerator.v:3502" *)
  wire _T_47;
  (* src = "crypto_accelerator.v:3716" *)
  wire _T_470;
  (* src = "crypto_accelerator.v:6083" *)
  wire [63:0] _T_4717;
  (* src = "crypto_accelerator.v:3717" *)
  wire _T_472;
  (* src = "crypto_accelerator.v:6084" *)
  wire [127:0] _T_4725;
  (* src = "crypto_accelerator.v:6085" *)
  wire [127:0] _T_4726;
  (* src = "crypto_accelerator.v:3718" *)
  wire _T_474;
  (* src = "crypto_accelerator.v:6102" *)
  wire _T_4747;
  (* src = "crypto_accelerator.v:3719" *)
  wire _T_476;
  wire [3:0] _T_4769;
  (* src = "crypto_accelerator.v:6104" *)
  wire _T_4770;
  (* src = "crypto_accelerator.v:6105" *)
  wire _T_4771;
  (* src = "crypto_accelerator.v:6108" *)
  wire _T_4775;
  (* src = "crypto_accelerator.v:6111" *)
  wire [5:0] _T_4778;
  (* src = "crypto_accelerator.v:3720" *)
  wire _T_478;
  (* src = "crypto_accelerator.v:3721" *)
  wire _T_480;
  (* src = "crypto_accelerator.v:3722" *)
  wire _T_482;
  (* src = "crypto_accelerator.v:3723" *)
  wire _T_484;
  (* src = "crypto_accelerator.v:3724" *)
  wire _T_486;
  (* src = "crypto_accelerator.v:3725" *)
  wire _T_488;
  (* src = "crypto_accelerator.v:3503" *)
  wire _T_49;
  (* src = "crypto_accelerator.v:3726" *)
  wire _T_490;
  (* src = "crypto_accelerator.v:3727" *)
  wire _T_492;
  (* src = "crypto_accelerator.v:3728" *)
  wire _T_494;
  (* src = "crypto_accelerator.v:3729" *)
  wire _T_496;
  (* src = "crypto_accelerator.v:3730" *)
  wire _T_498;
  (* src = "crypto_accelerator.v:3731" *)
  wire _T_500;
  (* src = "crypto_accelerator.v:3732" *)
  wire _T_502;
  (* src = "crypto_accelerator.v:3733" *)
  wire _T_504;
  (* src = "crypto_accelerator.v:3734" *)
  wire _T_506;
  (* src = "crypto_accelerator.v:3735" *)
  wire _T_508;
  (* src = "crypto_accelerator.v:3504" *)
  wire _T_51;
  (* src = "crypto_accelerator.v:3736" *)
  wire _T_510;
  (* src = "crypto_accelerator.v:3737" *)
  wire _T_512;
  (* src = "crypto_accelerator.v:3738" *)
  wire _T_514;
  (* src = "crypto_accelerator.v:3739" *)
  wire _T_516;
  (* src = "crypto_accelerator.v:3740" *)
  wire _T_518;
  (* src = "crypto_accelerator.v:3505" *)
  wire _T_52;
  (* src = "crypto_accelerator.v:3741" *)
  wire _T_520;
  (* src = "crypto_accelerator.v:3742" *)
  wire _T_522;
  (* src = "crypto_accelerator.v:3743" *)
  wire _T_524;
  (* src = "crypto_accelerator.v:3744" *)
  wire _T_526;
  (* src = "crypto_accelerator.v:3745" *)
  wire _T_528;
  (* src = "crypto_accelerator.v:3746" *)
  wire _T_530;
  (* src = "crypto_accelerator.v:3747" *)
  wire _T_532;
  (* src = "crypto_accelerator.v:3748" *)
  wire _T_534;
  (* src = "crypto_accelerator.v:3749" *)
  wire _T_536;
  (* src = "crypto_accelerator.v:3750" *)
  wire _T_538;
  (* src = "crypto_accelerator.v:3506" *)
  wire _T_54;
  (* src = "crypto_accelerator.v:3751" *)
  wire _T_540;
  (* src = "crypto_accelerator.v:3752" *)
  wire _T_542;
  (* src = "crypto_accelerator.v:3753" *)
  wire _T_544;
  (* src = "crypto_accelerator.v:3754" *)
  wire _T_546;
  (* src = "crypto_accelerator.v:3755" *)
  wire _T_548;
  (* src = "crypto_accelerator.v:3756" *)
  wire _T_550;
  (* src = "crypto_accelerator.v:3757" *)
  wire _T_552;
  (* src = "crypto_accelerator.v:3758" *)
  wire _T_554;
  (* src = "crypto_accelerator.v:3759" *)
  wire _T_556;
  (* src = "crypto_accelerator.v:3760" *)
  wire _T_558;
  (* src = "crypto_accelerator.v:3507" *)
  wire _T_56;
  (* src = "crypto_accelerator.v:3761" *)
  wire _T_560;
  (* src = "crypto_accelerator.v:3762" *)
  wire _T_562;
  (* src = "crypto_accelerator.v:3763" *)
  wire _T_564;
  (* src = "crypto_accelerator.v:3764" *)
  wire _T_566;
  (* src = "crypto_accelerator.v:3765" *)
  wire _T_567;
  (* src = "crypto_accelerator.v:3766" *)
  wire _T_568;
  (* src = "crypto_accelerator.v:3767" *)
  wire _T_569;
  (* src = "crypto_accelerator.v:3508" *)
  wire _T_57;
  (* src = "crypto_accelerator.v:3768" *)
  wire _T_570;
  (* src = "crypto_accelerator.v:3769" *)
  wire _T_571;
  (* src = "crypto_accelerator.v:3770" *)
  wire _T_572;
  (* src = "crypto_accelerator.v:3771" *)
  wire _T_573;
  (* src = "crypto_accelerator.v:3772" *)
  wire _T_574;
  (* src = "crypto_accelerator.v:3509" *)
  wire _T_59;
  (* src = "crypto_accelerator.v:3774" *)
  wire _T_599;
  (* src = "crypto_accelerator.v:3775" *)
  wire _T_601;
  (* src = "crypto_accelerator.v:3776" *)
  wire _T_602;
  (* src = "crypto_accelerator.v:3777" *)
  wire _T_604;
  (* src = "crypto_accelerator.v:3778" *)
  wire _T_605;
  (* src = "crypto_accelerator.v:3779" *)
  wire _T_607;
  (* src = "crypto_accelerator.v:3780" *)
  wire _T_609;
  (* src = "crypto_accelerator.v:3510" *)
  wire _T_61;
  (* src = "crypto_accelerator.v:3781" *)
  wire _T_610;
  (* src = "crypto_accelerator.v:3782" *)
  wire _T_612;
  (* src = "crypto_accelerator.v:3783" *)
  wire _T_614;
  (* src = "crypto_accelerator.v:3784" *)
  wire _T_615;
  (* src = "crypto_accelerator.v:3785" *)
  wire _T_617;
  (* src = "crypto_accelerator.v:3786" *)
  wire _T_619;
  (* src = "crypto_accelerator.v:3511" *)
  wire _T_62;
  (* src = "crypto_accelerator.v:3787" *)
  wire _T_620;
  (* src = "crypto_accelerator.v:3788" *)
  wire _T_622;
  (* src = "crypto_accelerator.v:3789" *)
  wire _T_624;
  (* src = "crypto_accelerator.v:3790" *)
  wire _T_626;
  (* src = "crypto_accelerator.v:3791" *)
  wire _T_628;
  (* src = "crypto_accelerator.v:3792" *)
  wire _T_629;
  (* src = "crypto_accelerator.v:3793" *)
  wire _T_631;
  (* src = "crypto_accelerator.v:3794" *)
  wire _T_633;
  (* src = "crypto_accelerator.v:3795" *)
  wire _T_634;
  (* src = "crypto_accelerator.v:3796" *)
  wire _T_636;
  (* src = "crypto_accelerator.v:3797" *)
  wire _T_638;
  (* src = "crypto_accelerator.v:3512" *)
  wire _T_64;
  (* src = "crypto_accelerator.v:3798" *)
  wire _T_640;
  (* src = "crypto_accelerator.v:3799" *)
  wire _T_641;
  (* src = "crypto_accelerator.v:3800" *)
  wire _T_643;
  (* src = "crypto_accelerator.v:3801" *)
  wire _T_644;
  (* src = "crypto_accelerator.v:3802" *)
  wire _T_646;
  (* src = "crypto_accelerator.v:3803" *)
  wire _T_647;
  (* src = "crypto_accelerator.v:3804" *)
  wire _T_649;
  (* src = "crypto_accelerator.v:3805" *)
  wire _T_651;
  (* src = "crypto_accelerator.v:3806" *)
  wire _T_653;
  (* src = "crypto_accelerator.v:3807" *)
  wire _T_655;
  (* src = "crypto_accelerator.v:3808" *)
  wire _T_657;
  (* src = "crypto_accelerator.v:3809" *)
  wire _T_659;
  (* src = "crypto_accelerator.v:3513" *)
  wire _T_66;
  (* src = "crypto_accelerator.v:3810" *)
  wire _T_661;
  (* src = "crypto_accelerator.v:3811" *)
  wire _T_663;
  (* src = "crypto_accelerator.v:3812" *)
  wire _T_665;
  (* src = "crypto_accelerator.v:3813" *)
  wire _T_667;
  (* src = "crypto_accelerator.v:3814" *)
  wire _T_669;
  (* src = "crypto_accelerator.v:3815" *)
  wire _T_671;
  (* src = "crypto_accelerator.v:3816" *)
  wire _T_673;
  (* src = "crypto_accelerator.v:3817" *)
  wire _T_675;
  (* src = "crypto_accelerator.v:3818" *)
  wire _T_677;
  (* src = "crypto_accelerator.v:3819" *)
  wire _T_679;
  (* src = "crypto_accelerator.v:3514" *)
  wire _T_68;
  (* src = "crypto_accelerator.v:3820" *)
  wire _T_681;
  (* src = "crypto_accelerator.v:3821" *)
  wire _T_683;
  (* src = "crypto_accelerator.v:3822" *)
  wire _T_685;
  (* src = "crypto_accelerator.v:3823" *)
  wire _T_687;
  (* src = "crypto_accelerator.v:3824" *)
  wire _T_689;
  (* src = "crypto_accelerator.v:3825" *)
  wire _T_691;
  (* src = "crypto_accelerator.v:3826" *)
  wire _T_693;
  (* src = "crypto_accelerator.v:3827" *)
  wire _T_695;
  (* src = "crypto_accelerator.v:3828" *)
  wire _T_697;
  (* src = "crypto_accelerator.v:3829" *)
  wire _T_699;
  (* src = "crypto_accelerator.v:3515" *)
  wire _T_70;
  (* src = "crypto_accelerator.v:3830" *)
  wire _T_701;
  (* src = "crypto_accelerator.v:3831" *)
  wire _T_703;
  (* src = "crypto_accelerator.v:3832" *)
  wire _T_705;
  (* src = "crypto_accelerator.v:3833" *)
  wire _T_707;
  (* src = "crypto_accelerator.v:3834" *)
  wire _T_709;
  (* src = "crypto_accelerator.v:3516" *)
  wire _T_71;
  (* src = "crypto_accelerator.v:3835" *)
  wire _T_711;
  (* src = "crypto_accelerator.v:3836" *)
  wire _T_713;
  (* src = "crypto_accelerator.v:3837" *)
  wire _T_715;
  (* src = "crypto_accelerator.v:3838" *)
  wire _T_717;
  (* src = "crypto_accelerator.v:3839" *)
  wire _T_719;
  (* src = "crypto_accelerator.v:3840" *)
  wire _T_721;
  (* src = "crypto_accelerator.v:3841" *)
  wire _T_723;
  (* src = "crypto_accelerator.v:3842" *)
  wire _T_725;
  (* src = "crypto_accelerator.v:3843" *)
  wire _T_727;
  (* src = "crypto_accelerator.v:3844" *)
  wire _T_729;
  (* src = "crypto_accelerator.v:3517" *)
  wire _T_73;
  (* src = "crypto_accelerator.v:3845" *)
  wire _T_731;
  (* src = "crypto_accelerator.v:3846" *)
  wire _T_733;
  (* src = "crypto_accelerator.v:3847" *)
  wire _T_735;
  (* src = "crypto_accelerator.v:3848" *)
  wire _T_737;
  (* src = "crypto_accelerator.v:3849" *)
  wire _T_739;
  (* src = "crypto_accelerator.v:3850" *)
  wire _T_741;
  (* src = "crypto_accelerator.v:3851" *)
  wire _T_743;
  (* src = "crypto_accelerator.v:3852" *)
  wire _T_745;
  (* src = "crypto_accelerator.v:3853" *)
  wire _T_747;
  (* src = "crypto_accelerator.v:3854" *)
  wire _T_749;
  (* src = "crypto_accelerator.v:3518" *)
  wire _T_75;
  (* src = "crypto_accelerator.v:3855" *)
  wire _T_751;
  (* src = "crypto_accelerator.v:3856" *)
  wire _T_753;
  (* src = "crypto_accelerator.v:3857" *)
  wire _T_755;
  (* src = "crypto_accelerator.v:3858" *)
  wire _T_757;
  (* src = "crypto_accelerator.v:3859" *)
  wire _T_759;
  (* src = "crypto_accelerator.v:3519" *)
  wire _T_76;
  (* src = "crypto_accelerator.v:3860" *)
  wire _T_761;
  (* src = "crypto_accelerator.v:3861" *)
  wire _T_763;
  (* src = "crypto_accelerator.v:3862" *)
  wire _T_765;
  (* src = "crypto_accelerator.v:3863" *)
  wire _T_767;
  (* src = "crypto_accelerator.v:3864" *)
  wire _T_769;
  (* src = "crypto_accelerator.v:3865" *)
  wire _T_771;
  (* src = "crypto_accelerator.v:3866" *)
  wire _T_773;
  (* src = "crypto_accelerator.v:3867" *)
  wire _T_775;
  (* src = "crypto_accelerator.v:3868" *)
  wire _T_777;
  (* src = "crypto_accelerator.v:3869" *)
  wire _T_779;
  (* src = "crypto_accelerator.v:3520" *)
  wire _T_78;
  (* src = "crypto_accelerator.v:3870" *)
  wire _T_781;
  (* src = "crypto_accelerator.v:3871" *)
  wire _T_783;
  (* src = "crypto_accelerator.v:3872" *)
  wire _T_785;
  (* src = "crypto_accelerator.v:3873" *)
  wire _T_787;
  (* src = "crypto_accelerator.v:3874" *)
  wire _T_789;
  (* src = "crypto_accelerator.v:3875" *)
  wire _T_791;
  (* src = "crypto_accelerator.v:3876" *)
  wire _T_793;
  (* src = "crypto_accelerator.v:3877" *)
  wire _T_795;
  (* src = "crypto_accelerator.v:3878" *)
  wire _T_797;
  (* src = "crypto_accelerator.v:3879" *)
  wire _T_799;
  (* src = "crypto_accelerator.v:3521" *)
  wire _T_80;
  (* src = "crypto_accelerator.v:3880" *)
  wire _T_801;
  (* src = "crypto_accelerator.v:3881" *)
  wire _T_803;
  (* src = "crypto_accelerator.v:3882" *)
  wire _T_805;
  (* src = "crypto_accelerator.v:3883" *)
  wire _T_807;
  (* src = "crypto_accelerator.v:3884" *)
  wire _T_809;
  (* src = "crypto_accelerator.v:3885" *)
  wire _T_811;
  (* src = "crypto_accelerator.v:3886" *)
  wire _T_813;
  (* src = "crypto_accelerator.v:3887" *)
  wire _T_815;
  (* src = "crypto_accelerator.v:3888" *)
  wire _T_817;
  (* src = "crypto_accelerator.v:3889" *)
  wire _T_819;
  (* src = "crypto_accelerator.v:3522" *)
  wire _T_82;
  (* src = "crypto_accelerator.v:3890" *)
  wire _T_821;
  (* src = "crypto_accelerator.v:3891" *)
  wire _T_823;
  (* src = "crypto_accelerator.v:3892" *)
  wire _T_825;
  (* src = "crypto_accelerator.v:3893" *)
  wire _T_827;
  (* src = "crypto_accelerator.v:3894" *)
  wire _T_829;
  (* src = "crypto_accelerator.v:3523" *)
  wire _T_83;
  (* src = "crypto_accelerator.v:3895" *)
  wire _T_831;
  (* src = "crypto_accelerator.v:3896" *)
  wire _T_833;
  (* src = "crypto_accelerator.v:3897" *)
  wire _T_835;
  (* src = "crypto_accelerator.v:3898" *)
  wire _T_837;
  (* src = "crypto_accelerator.v:3899" *)
  wire _T_839;
  (* src = "crypto_accelerator.v:3900" *)
  wire _T_841;
  (* src = "crypto_accelerator.v:3901" *)
  wire _T_843;
  (* src = "crypto_accelerator.v:3902" *)
  wire _T_845;
  (* src = "crypto_accelerator.v:3903" *)
  wire _T_846;
  (* src = "crypto_accelerator.v:3904" *)
  wire _T_847;
  (* src = "crypto_accelerator.v:3905" *)
  wire _T_848;
  (* src = "crypto_accelerator.v:3906" *)
  wire _T_849;
  (* src = "crypto_accelerator.v:3524" *)
  wire _T_85;
  (* src = "crypto_accelerator.v:3907" *)
  wire _T_850;
  (* src = "crypto_accelerator.v:3908" *)
  wire _T_851;
  (* src = "crypto_accelerator.v:3909" *)
  wire _T_852;
  (* src = "crypto_accelerator.v:3910" *)
  wire _T_853;
  (* src = "crypto_accelerator.v:3525" *)
  wire _T_86;
  (* src = "crypto_accelerator.v:3912" *)
  wire _T_878;
  (* src = "crypto_accelerator.v:3526" *)
  wire _T_88;
  (* src = "crypto_accelerator.v:3913" *)
  wire _T_880;
  (* src = "crypto_accelerator.v:3914" *)
  wire _T_881;
  (* src = "crypto_accelerator.v:3915" *)
  wire _T_883;
  (* src = "crypto_accelerator.v:3916" *)
  wire _T_884;
  (* src = "crypto_accelerator.v:3917" *)
  wire _T_886;
  (* src = "crypto_accelerator.v:3918" *)
  wire _T_888;
  (* src = "crypto_accelerator.v:3919" *)
  wire _T_889;
  (* src = "crypto_accelerator.v:3527" *)
  wire _T_89;
  (* src = "crypto_accelerator.v:3920" *)
  wire _T_891;
  (* src = "crypto_accelerator.v:3921" *)
  wire _T_893;
  (* src = "crypto_accelerator.v:3922" *)
  wire _T_894;
  (* src = "crypto_accelerator.v:3923" *)
  wire _T_896;
  (* src = "crypto_accelerator.v:3924" *)
  wire _T_898;
  (* src = "crypto_accelerator.v:3925" *)
  wire _T_899;
  (* src = "crypto_accelerator.v:3926" *)
  wire _T_901;
  (* src = "crypto_accelerator.v:3927" *)
  wire _T_903;
  (* src = "crypto_accelerator.v:3928" *)
  wire _T_905;
  (* src = "crypto_accelerator.v:3929" *)
  wire _T_907;
  (* src = "crypto_accelerator.v:3930" *)
  wire _T_908;
  (* src = "crypto_accelerator.v:3528" *)
  wire _T_91;
  (* src = "crypto_accelerator.v:3931" *)
  wire _T_910;
  (* src = "crypto_accelerator.v:3932" *)
  wire _T_912;
  (* src = "crypto_accelerator.v:3933" *)
  wire _T_913;
  (* src = "crypto_accelerator.v:3934" *)
  wire _T_915;
  (* src = "crypto_accelerator.v:3935" *)
  wire _T_917;
  (* src = "crypto_accelerator.v:3936" *)
  wire _T_919;
  (* src = "crypto_accelerator.v:3937" *)
  wire _T_920;
  (* src = "crypto_accelerator.v:3938" *)
  wire _T_922;
  (* src = "crypto_accelerator.v:3939" *)
  wire _T_923;
  (* src = "crypto_accelerator.v:3940" *)
  wire _T_925;
  (* src = "crypto_accelerator.v:3941" *)
  wire _T_926;
  (* src = "crypto_accelerator.v:3942" *)
  wire _T_928;
  (* src = "crypto_accelerator.v:3529" *)
  wire _T_93;
  (* src = "crypto_accelerator.v:3943" *)
  wire _T_930;
  (* src = "crypto_accelerator.v:3944" *)
  wire _T_932;
  (* src = "crypto_accelerator.v:3945" *)
  wire _T_934;
  (* src = "crypto_accelerator.v:3946" *)
  wire _T_936;
  (* src = "crypto_accelerator.v:3947" *)
  wire _T_938;
  (* src = "crypto_accelerator.v:3948" *)
  wire _T_940;
  (* src = "crypto_accelerator.v:3949" *)
  wire _T_942;
  (* src = "crypto_accelerator.v:3950" *)
  wire _T_944;
  (* src = "crypto_accelerator.v:3951" *)
  wire _T_946;
  (* src = "crypto_accelerator.v:3952" *)
  wire _T_948;
  (* src = "crypto_accelerator.v:3530" *)
  wire _T_95;
  (* src = "crypto_accelerator.v:3953" *)
  wire _T_950;
  (* src = "crypto_accelerator.v:3954" *)
  wire _T_952;
  (* src = "crypto_accelerator.v:3955" *)
  wire _T_954;
  (* src = "crypto_accelerator.v:3956" *)
  wire _T_956;
  (* src = "crypto_accelerator.v:3957" *)
  wire _T_958;
  (* src = "crypto_accelerator.v:3958" *)
  wire _T_960;
  (* src = "crypto_accelerator.v:3959" *)
  wire _T_962;
  (* src = "crypto_accelerator.v:3960" *)
  wire _T_964;
  (* src = "crypto_accelerator.v:3961" *)
  wire _T_966;
  (* src = "crypto_accelerator.v:3962" *)
  wire _T_968;
  (* src = "crypto_accelerator.v:3531" *)
  wire _T_97;
  (* src = "crypto_accelerator.v:3963" *)
  wire _T_970;
  (* src = "crypto_accelerator.v:3964" *)
  wire _T_972;
  (* src = "crypto_accelerator.v:3965" *)
  wire _T_974;
  (* src = "crypto_accelerator.v:3966" *)
  wire _T_976;
  (* src = "crypto_accelerator.v:3967" *)
  wire _T_978;
  (* src = "crypto_accelerator.v:3968" *)
  wire _T_980;
  (* src = "crypto_accelerator.v:3969" *)
  wire _T_982;
  (* src = "crypto_accelerator.v:3970" *)
  wire _T_984;
  (* src = "crypto_accelerator.v:3971" *)
  wire _T_986;
  (* src = "crypto_accelerator.v:3972" *)
  wire _T_988;
  (* src = "crypto_accelerator.v:3532" *)
  wire _T_99;
  (* src = "crypto_accelerator.v:3973" *)
  wire _T_990;
  (* src = "crypto_accelerator.v:3974" *)
  wire _T_992;
  (* src = "crypto_accelerator.v:3975" *)
  wire _T_994;
  (* src = "crypto_accelerator.v:3976" *)
  wire _T_996;
  (* src = "crypto_accelerator.v:3977" *)
  wire _T_998;
  (* src = "crypto_accelerator.v:3170" *)
  input clock;
  (* src = "crypto_accelerator.v:3479" *)
  reg [127:0] ctSaved;
  (* src = "crypto_accelerator.v:6086" *)
  wire [7:0] finalOut_0_0;
  (* src = "crypto_accelerator.v:6087" *)
  wire [7:0] finalOut_0_1;
  (* src = "crypto_accelerator.v:6088" *)
  wire [7:0] finalOut_0_2;
  (* src = "crypto_accelerator.v:6089" *)
  wire [7:0] finalOut_0_3;
  (* src = "crypto_accelerator.v:6090" *)
  wire [7:0] finalOut_1_0;
  (* src = "crypto_accelerator.v:6091" *)
  wire [7:0] finalOut_1_1;
  (* src = "crypto_accelerator.v:6092" *)
  wire [7:0] finalOut_1_2;
  (* src = "crypto_accelerator.v:6093" *)
  wire [7:0] finalOut_1_3;
  (* src = "crypto_accelerator.v:6094" *)
  wire [7:0] finalOut_2_0;
  (* src = "crypto_accelerator.v:6095" *)
  wire [7:0] finalOut_2_1;
  (* src = "crypto_accelerator.v:6096" *)
  wire [7:0] finalOut_2_2;
  (* src = "crypto_accelerator.v:6097" *)
  wire [7:0] finalOut_2_3;
  (* src = "crypto_accelerator.v:6098" *)
  wire [7:0] finalOut_3_0;
  (* src = "crypto_accelerator.v:6099" *)
  wire [7:0] finalOut_3_1;
  (* src = "crypto_accelerator.v:6100" *)
  wire [7:0] finalOut_3_2;
  (* src = "crypto_accelerator.v:6101" *)
  wire [7:0] finalOut_3_3;
  (* src = "crypto_accelerator.v:3415" *)
  input io_aes256;
  (* src = "crypto_accelerator.v:3172" *)
  input [127:0] io_dataIn;
  (* src = "crypto_accelerator.v:3420" *)
  output [127:0] io_dataOut;
  (* src = "crypto_accelerator.v:3174" *)
  input io_dataValid;
  (* src = "crypto_accelerator.v:3173" *)
  input [127:0] io_ivIn;
  (* src = "crypto_accelerator.v:3421" *)
  output [127:0] io_ivOut;
  (* src = "crypto_accelerator.v:3175" *)
  input [7:0] io_keys_0_0_0;
  (* src = "crypto_accelerator.v:3176" *)
  input [7:0] io_keys_0_0_1;
  (* src = "crypto_accelerator.v:3177" *)
  input [7:0] io_keys_0_0_2;
  (* src = "crypto_accelerator.v:3178" *)
  input [7:0] io_keys_0_0_3;
  (* src = "crypto_accelerator.v:3179" *)
  input [7:0] io_keys_0_1_0;
  (* src = "crypto_accelerator.v:3180" *)
  input [7:0] io_keys_0_1_1;
  (* src = "crypto_accelerator.v:3181" *)
  input [7:0] io_keys_0_1_2;
  (* src = "crypto_accelerator.v:3182" *)
  input [7:0] io_keys_0_1_3;
  (* src = "crypto_accelerator.v:3183" *)
  input [7:0] io_keys_0_2_0;
  (* src = "crypto_accelerator.v:3184" *)
  input [7:0] io_keys_0_2_1;
  (* src = "crypto_accelerator.v:3185" *)
  input [7:0] io_keys_0_2_2;
  (* src = "crypto_accelerator.v:3186" *)
  input [7:0] io_keys_0_2_3;
  (* src = "crypto_accelerator.v:3187" *)
  input [7:0] io_keys_0_3_0;
  (* src = "crypto_accelerator.v:3188" *)
  input [7:0] io_keys_0_3_1;
  (* src = "crypto_accelerator.v:3189" *)
  input [7:0] io_keys_0_3_2;
  (* src = "crypto_accelerator.v:3190" *)
  input [7:0] io_keys_0_3_3;
  (* src = "crypto_accelerator.v:3335" *)
  input [7:0] io_keys_10_0_0;
  (* src = "crypto_accelerator.v:3336" *)
  input [7:0] io_keys_10_0_1;
  (* src = "crypto_accelerator.v:3337" *)
  input [7:0] io_keys_10_0_2;
  (* src = "crypto_accelerator.v:3338" *)
  input [7:0] io_keys_10_0_3;
  (* src = "crypto_accelerator.v:3339" *)
  input [7:0] io_keys_10_1_0;
  (* src = "crypto_accelerator.v:3340" *)
  input [7:0] io_keys_10_1_1;
  (* src = "crypto_accelerator.v:3341" *)
  input [7:0] io_keys_10_1_2;
  (* src = "crypto_accelerator.v:3342" *)
  input [7:0] io_keys_10_1_3;
  (* src = "crypto_accelerator.v:3343" *)
  input [7:0] io_keys_10_2_0;
  (* src = "crypto_accelerator.v:3344" *)
  input [7:0] io_keys_10_2_1;
  (* src = "crypto_accelerator.v:3345" *)
  input [7:0] io_keys_10_2_2;
  (* src = "crypto_accelerator.v:3346" *)
  input [7:0] io_keys_10_2_3;
  (* src = "crypto_accelerator.v:3347" *)
  input [7:0] io_keys_10_3_0;
  (* src = "crypto_accelerator.v:3348" *)
  input [7:0] io_keys_10_3_1;
  (* src = "crypto_accelerator.v:3349" *)
  input [7:0] io_keys_10_3_2;
  (* src = "crypto_accelerator.v:3350" *)
  input [7:0] io_keys_10_3_3;
  (* src = "crypto_accelerator.v:3351" *)
  input [7:0] io_keys_11_0_0;
  (* src = "crypto_accelerator.v:3352" *)
  input [7:0] io_keys_11_0_1;
  (* src = "crypto_accelerator.v:3353" *)
  input [7:0] io_keys_11_0_2;
  (* src = "crypto_accelerator.v:3354" *)
  input [7:0] io_keys_11_0_3;
  (* src = "crypto_accelerator.v:3355" *)
  input [7:0] io_keys_11_1_0;
  (* src = "crypto_accelerator.v:3356" *)
  input [7:0] io_keys_11_1_1;
  (* src = "crypto_accelerator.v:3357" *)
  input [7:0] io_keys_11_1_2;
  (* src = "crypto_accelerator.v:3358" *)
  input [7:0] io_keys_11_1_3;
  (* src = "crypto_accelerator.v:3359" *)
  input [7:0] io_keys_11_2_0;
  (* src = "crypto_accelerator.v:3360" *)
  input [7:0] io_keys_11_2_1;
  (* src = "crypto_accelerator.v:3361" *)
  input [7:0] io_keys_11_2_2;
  (* src = "crypto_accelerator.v:3362" *)
  input [7:0] io_keys_11_2_3;
  (* src = "crypto_accelerator.v:3363" *)
  input [7:0] io_keys_11_3_0;
  (* src = "crypto_accelerator.v:3364" *)
  input [7:0] io_keys_11_3_1;
  (* src = "crypto_accelerator.v:3365" *)
  input [7:0] io_keys_11_3_2;
  (* src = "crypto_accelerator.v:3366" *)
  input [7:0] io_keys_11_3_3;
  (* src = "crypto_accelerator.v:3367" *)
  input [7:0] io_keys_12_0_0;
  (* src = "crypto_accelerator.v:3368" *)
  input [7:0] io_keys_12_0_1;
  (* src = "crypto_accelerator.v:3369" *)
  input [7:0] io_keys_12_0_2;
  (* src = "crypto_accelerator.v:3370" *)
  input [7:0] io_keys_12_0_3;
  (* src = "crypto_accelerator.v:3371" *)
  input [7:0] io_keys_12_1_0;
  (* src = "crypto_accelerator.v:3372" *)
  input [7:0] io_keys_12_1_1;
  (* src = "crypto_accelerator.v:3373" *)
  input [7:0] io_keys_12_1_2;
  (* src = "crypto_accelerator.v:3374" *)
  input [7:0] io_keys_12_1_3;
  (* src = "crypto_accelerator.v:3375" *)
  input [7:0] io_keys_12_2_0;
  (* src = "crypto_accelerator.v:3376" *)
  input [7:0] io_keys_12_2_1;
  (* src = "crypto_accelerator.v:3377" *)
  input [7:0] io_keys_12_2_2;
  (* src = "crypto_accelerator.v:3378" *)
  input [7:0] io_keys_12_2_3;
  (* src = "crypto_accelerator.v:3379" *)
  input [7:0] io_keys_12_3_0;
  (* src = "crypto_accelerator.v:3380" *)
  input [7:0] io_keys_12_3_1;
  (* src = "crypto_accelerator.v:3381" *)
  input [7:0] io_keys_12_3_2;
  (* src = "crypto_accelerator.v:3382" *)
  input [7:0] io_keys_12_3_3;
  (* src = "crypto_accelerator.v:3383" *)
  input [7:0] io_keys_13_0_0;
  (* src = "crypto_accelerator.v:3384" *)
  input [7:0] io_keys_13_0_1;
  (* src = "crypto_accelerator.v:3385" *)
  input [7:0] io_keys_13_0_2;
  (* src = "crypto_accelerator.v:3386" *)
  input [7:0] io_keys_13_0_3;
  (* src = "crypto_accelerator.v:3387" *)
  input [7:0] io_keys_13_1_0;
  (* src = "crypto_accelerator.v:3388" *)
  input [7:0] io_keys_13_1_1;
  (* src = "crypto_accelerator.v:3389" *)
  input [7:0] io_keys_13_1_2;
  (* src = "crypto_accelerator.v:3390" *)
  input [7:0] io_keys_13_1_3;
  (* src = "crypto_accelerator.v:3391" *)
  input [7:0] io_keys_13_2_0;
  (* src = "crypto_accelerator.v:3392" *)
  input [7:0] io_keys_13_2_1;
  (* src = "crypto_accelerator.v:3393" *)
  input [7:0] io_keys_13_2_2;
  (* src = "crypto_accelerator.v:3394" *)
  input [7:0] io_keys_13_2_3;
  (* src = "crypto_accelerator.v:3395" *)
  input [7:0] io_keys_13_3_0;
  (* src = "crypto_accelerator.v:3396" *)
  input [7:0] io_keys_13_3_1;
  (* src = "crypto_accelerator.v:3397" *)
  input [7:0] io_keys_13_3_2;
  (* src = "crypto_accelerator.v:3398" *)
  input [7:0] io_keys_13_3_3;
  (* src = "crypto_accelerator.v:3399" *)
  input [7:0] io_keys_14_0_0;
  (* src = "crypto_accelerator.v:3400" *)
  input [7:0] io_keys_14_0_1;
  (* src = "crypto_accelerator.v:3401" *)
  input [7:0] io_keys_14_0_2;
  (* src = "crypto_accelerator.v:3402" *)
  input [7:0] io_keys_14_0_3;
  (* src = "crypto_accelerator.v:3403" *)
  input [7:0] io_keys_14_1_0;
  (* src = "crypto_accelerator.v:3404" *)
  input [7:0] io_keys_14_1_1;
  (* src = "crypto_accelerator.v:3405" *)
  input [7:0] io_keys_14_1_2;
  (* src = "crypto_accelerator.v:3406" *)
  input [7:0] io_keys_14_1_3;
  (* src = "crypto_accelerator.v:3407" *)
  input [7:0] io_keys_14_2_0;
  (* src = "crypto_accelerator.v:3408" *)
  input [7:0] io_keys_14_2_1;
  (* src = "crypto_accelerator.v:3409" *)
  input [7:0] io_keys_14_2_2;
  (* src = "crypto_accelerator.v:3410" *)
  input [7:0] io_keys_14_2_3;
  (* src = "crypto_accelerator.v:3411" *)
  input [7:0] io_keys_14_3_0;
  (* src = "crypto_accelerator.v:3412" *)
  input [7:0] io_keys_14_3_1;
  (* src = "crypto_accelerator.v:3413" *)
  input [7:0] io_keys_14_3_2;
  (* src = "crypto_accelerator.v:3414" *)
  input [7:0] io_keys_14_3_3;
  (* src = "crypto_accelerator.v:3191" *)
  input [7:0] io_keys_1_0_0;
  (* src = "crypto_accelerator.v:3192" *)
  input [7:0] io_keys_1_0_1;
  (* src = "crypto_accelerator.v:3193" *)
  input [7:0] io_keys_1_0_2;
  (* src = "crypto_accelerator.v:3194" *)
  input [7:0] io_keys_1_0_3;
  (* src = "crypto_accelerator.v:3195" *)
  input [7:0] io_keys_1_1_0;
  (* src = "crypto_accelerator.v:3196" *)
  input [7:0] io_keys_1_1_1;
  (* src = "crypto_accelerator.v:3197" *)
  input [7:0] io_keys_1_1_2;
  (* src = "crypto_accelerator.v:3198" *)
  input [7:0] io_keys_1_1_3;
  (* src = "crypto_accelerator.v:3199" *)
  input [7:0] io_keys_1_2_0;
  (* src = "crypto_accelerator.v:3200" *)
  input [7:0] io_keys_1_2_1;
  (* src = "crypto_accelerator.v:3201" *)
  input [7:0] io_keys_1_2_2;
  (* src = "crypto_accelerator.v:3202" *)
  input [7:0] io_keys_1_2_3;
  (* src = "crypto_accelerator.v:3203" *)
  input [7:0] io_keys_1_3_0;
  (* src = "crypto_accelerator.v:3204" *)
  input [7:0] io_keys_1_3_1;
  (* src = "crypto_accelerator.v:3205" *)
  input [7:0] io_keys_1_3_2;
  (* src = "crypto_accelerator.v:3206" *)
  input [7:0] io_keys_1_3_3;
  (* src = "crypto_accelerator.v:3207" *)
  input [7:0] io_keys_2_0_0;
  (* src = "crypto_accelerator.v:3208" *)
  input [7:0] io_keys_2_0_1;
  (* src = "crypto_accelerator.v:3209" *)
  input [7:0] io_keys_2_0_2;
  (* src = "crypto_accelerator.v:3210" *)
  input [7:0] io_keys_2_0_3;
  (* src = "crypto_accelerator.v:3211" *)
  input [7:0] io_keys_2_1_0;
  (* src = "crypto_accelerator.v:3212" *)
  input [7:0] io_keys_2_1_1;
  (* src = "crypto_accelerator.v:3213" *)
  input [7:0] io_keys_2_1_2;
  (* src = "crypto_accelerator.v:3214" *)
  input [7:0] io_keys_2_1_3;
  (* src = "crypto_accelerator.v:3215" *)
  input [7:0] io_keys_2_2_0;
  (* src = "crypto_accelerator.v:3216" *)
  input [7:0] io_keys_2_2_1;
  (* src = "crypto_accelerator.v:3217" *)
  input [7:0] io_keys_2_2_2;
  (* src = "crypto_accelerator.v:3218" *)
  input [7:0] io_keys_2_2_3;
  (* src = "crypto_accelerator.v:3219" *)
  input [7:0] io_keys_2_3_0;
  (* src = "crypto_accelerator.v:3220" *)
  input [7:0] io_keys_2_3_1;
  (* src = "crypto_accelerator.v:3221" *)
  input [7:0] io_keys_2_3_2;
  (* src = "crypto_accelerator.v:3222" *)
  input [7:0] io_keys_2_3_3;
  (* src = "crypto_accelerator.v:3223" *)
  input [7:0] io_keys_3_0_0;
  (* src = "crypto_accelerator.v:3224" *)
  input [7:0] io_keys_3_0_1;
  (* src = "crypto_accelerator.v:3225" *)
  input [7:0] io_keys_3_0_2;
  (* src = "crypto_accelerator.v:3226" *)
  input [7:0] io_keys_3_0_3;
  (* src = "crypto_accelerator.v:3227" *)
  input [7:0] io_keys_3_1_0;
  (* src = "crypto_accelerator.v:3228" *)
  input [7:0] io_keys_3_1_1;
  (* src = "crypto_accelerator.v:3229" *)
  input [7:0] io_keys_3_1_2;
  (* src = "crypto_accelerator.v:3230" *)
  input [7:0] io_keys_3_1_3;
  (* src = "crypto_accelerator.v:3231" *)
  input [7:0] io_keys_3_2_0;
  (* src = "crypto_accelerator.v:3232" *)
  input [7:0] io_keys_3_2_1;
  (* src = "crypto_accelerator.v:3233" *)
  input [7:0] io_keys_3_2_2;
  (* src = "crypto_accelerator.v:3234" *)
  input [7:0] io_keys_3_2_3;
  (* src = "crypto_accelerator.v:3235" *)
  input [7:0] io_keys_3_3_0;
  (* src = "crypto_accelerator.v:3236" *)
  input [7:0] io_keys_3_3_1;
  (* src = "crypto_accelerator.v:3237" *)
  input [7:0] io_keys_3_3_2;
  (* src = "crypto_accelerator.v:3238" *)
  input [7:0] io_keys_3_3_3;
  (* src = "crypto_accelerator.v:3239" *)
  input [7:0] io_keys_4_0_0;
  (* src = "crypto_accelerator.v:3240" *)
  input [7:0] io_keys_4_0_1;
  (* src = "crypto_accelerator.v:3241" *)
  input [7:0] io_keys_4_0_2;
  (* src = "crypto_accelerator.v:3242" *)
  input [7:0] io_keys_4_0_3;
  (* src = "crypto_accelerator.v:3243" *)
  input [7:0] io_keys_4_1_0;
  (* src = "crypto_accelerator.v:3244" *)
  input [7:0] io_keys_4_1_1;
  (* src = "crypto_accelerator.v:3245" *)
  input [7:0] io_keys_4_1_2;
  (* src = "crypto_accelerator.v:3246" *)
  input [7:0] io_keys_4_1_3;
  (* src = "crypto_accelerator.v:3247" *)
  input [7:0] io_keys_4_2_0;
  (* src = "crypto_accelerator.v:3248" *)
  input [7:0] io_keys_4_2_1;
  (* src = "crypto_accelerator.v:3249" *)
  input [7:0] io_keys_4_2_2;
  (* src = "crypto_accelerator.v:3250" *)
  input [7:0] io_keys_4_2_3;
  (* src = "crypto_accelerator.v:3251" *)
  input [7:0] io_keys_4_3_0;
  (* src = "crypto_accelerator.v:3252" *)
  input [7:0] io_keys_4_3_1;
  (* src = "crypto_accelerator.v:3253" *)
  input [7:0] io_keys_4_3_2;
  (* src = "crypto_accelerator.v:3254" *)
  input [7:0] io_keys_4_3_3;
  (* src = "crypto_accelerator.v:3255" *)
  input [7:0] io_keys_5_0_0;
  (* src = "crypto_accelerator.v:3256" *)
  input [7:0] io_keys_5_0_1;
  (* src = "crypto_accelerator.v:3257" *)
  input [7:0] io_keys_5_0_2;
  (* src = "crypto_accelerator.v:3258" *)
  input [7:0] io_keys_5_0_3;
  (* src = "crypto_accelerator.v:3259" *)
  input [7:0] io_keys_5_1_0;
  (* src = "crypto_accelerator.v:3260" *)
  input [7:0] io_keys_5_1_1;
  (* src = "crypto_accelerator.v:3261" *)
  input [7:0] io_keys_5_1_2;
  (* src = "crypto_accelerator.v:3262" *)
  input [7:0] io_keys_5_1_3;
  (* src = "crypto_accelerator.v:3263" *)
  input [7:0] io_keys_5_2_0;
  (* src = "crypto_accelerator.v:3264" *)
  input [7:0] io_keys_5_2_1;
  (* src = "crypto_accelerator.v:3265" *)
  input [7:0] io_keys_5_2_2;
  (* src = "crypto_accelerator.v:3266" *)
  input [7:0] io_keys_5_2_3;
  (* src = "crypto_accelerator.v:3267" *)
  input [7:0] io_keys_5_3_0;
  (* src = "crypto_accelerator.v:3268" *)
  input [7:0] io_keys_5_3_1;
  (* src = "crypto_accelerator.v:3269" *)
  input [7:0] io_keys_5_3_2;
  (* src = "crypto_accelerator.v:3270" *)
  input [7:0] io_keys_5_3_3;
  (* src = "crypto_accelerator.v:3271" *)
  input [7:0] io_keys_6_0_0;
  (* src = "crypto_accelerator.v:3272" *)
  input [7:0] io_keys_6_0_1;
  (* src = "crypto_accelerator.v:3273" *)
  input [7:0] io_keys_6_0_2;
  (* src = "crypto_accelerator.v:3274" *)
  input [7:0] io_keys_6_0_3;
  (* src = "crypto_accelerator.v:3275" *)
  input [7:0] io_keys_6_1_0;
  (* src = "crypto_accelerator.v:3276" *)
  input [7:0] io_keys_6_1_1;
  (* src = "crypto_accelerator.v:3277" *)
  input [7:0] io_keys_6_1_2;
  (* src = "crypto_accelerator.v:3278" *)
  input [7:0] io_keys_6_1_3;
  (* src = "crypto_accelerator.v:3279" *)
  input [7:0] io_keys_6_2_0;
  (* src = "crypto_accelerator.v:3280" *)
  input [7:0] io_keys_6_2_1;
  (* src = "crypto_accelerator.v:3281" *)
  input [7:0] io_keys_6_2_2;
  (* src = "crypto_accelerator.v:3282" *)
  input [7:0] io_keys_6_2_3;
  (* src = "crypto_accelerator.v:3283" *)
  input [7:0] io_keys_6_3_0;
  (* src = "crypto_accelerator.v:3284" *)
  input [7:0] io_keys_6_3_1;
  (* src = "crypto_accelerator.v:3285" *)
  input [7:0] io_keys_6_3_2;
  (* src = "crypto_accelerator.v:3286" *)
  input [7:0] io_keys_6_3_3;
  (* src = "crypto_accelerator.v:3287" *)
  input [7:0] io_keys_7_0_0;
  (* src = "crypto_accelerator.v:3288" *)
  input [7:0] io_keys_7_0_1;
  (* src = "crypto_accelerator.v:3289" *)
  input [7:0] io_keys_7_0_2;
  (* src = "crypto_accelerator.v:3290" *)
  input [7:0] io_keys_7_0_3;
  (* src = "crypto_accelerator.v:3291" *)
  input [7:0] io_keys_7_1_0;
  (* src = "crypto_accelerator.v:3292" *)
  input [7:0] io_keys_7_1_1;
  (* src = "crypto_accelerator.v:3293" *)
  input [7:0] io_keys_7_1_2;
  (* src = "crypto_accelerator.v:3294" *)
  input [7:0] io_keys_7_1_3;
  (* src = "crypto_accelerator.v:3295" *)
  input [7:0] io_keys_7_2_0;
  (* src = "crypto_accelerator.v:3296" *)
  input [7:0] io_keys_7_2_1;
  (* src = "crypto_accelerator.v:3297" *)
  input [7:0] io_keys_7_2_2;
  (* src = "crypto_accelerator.v:3298" *)
  input [7:0] io_keys_7_2_3;
  (* src = "crypto_accelerator.v:3299" *)
  input [7:0] io_keys_7_3_0;
  (* src = "crypto_accelerator.v:3300" *)
  input [7:0] io_keys_7_3_1;
  (* src = "crypto_accelerator.v:3301" *)
  input [7:0] io_keys_7_3_2;
  (* src = "crypto_accelerator.v:3302" *)
  input [7:0] io_keys_7_3_3;
  (* src = "crypto_accelerator.v:3303" *)
  input [7:0] io_keys_8_0_0;
  (* src = "crypto_accelerator.v:3304" *)
  input [7:0] io_keys_8_0_1;
  (* src = "crypto_accelerator.v:3305" *)
  input [7:0] io_keys_8_0_2;
  (* src = "crypto_accelerator.v:3306" *)
  input [7:0] io_keys_8_0_3;
  (* src = "crypto_accelerator.v:3307" *)
  input [7:0] io_keys_8_1_0;
  (* src = "crypto_accelerator.v:3308" *)
  input [7:0] io_keys_8_1_1;
  (* src = "crypto_accelerator.v:3309" *)
  input [7:0] io_keys_8_1_2;
  (* src = "crypto_accelerator.v:3310" *)
  input [7:0] io_keys_8_1_3;
  (* src = "crypto_accelerator.v:3311" *)
  input [7:0] io_keys_8_2_0;
  (* src = "crypto_accelerator.v:3312" *)
  input [7:0] io_keys_8_2_1;
  (* src = "crypto_accelerator.v:3313" *)
  input [7:0] io_keys_8_2_2;
  (* src = "crypto_accelerator.v:3314" *)
  input [7:0] io_keys_8_2_3;
  (* src = "crypto_accelerator.v:3315" *)
  input [7:0] io_keys_8_3_0;
  (* src = "crypto_accelerator.v:3316" *)
  input [7:0] io_keys_8_3_1;
  (* src = "crypto_accelerator.v:3317" *)
  input [7:0] io_keys_8_3_2;
  (* src = "crypto_accelerator.v:3318" *)
  input [7:0] io_keys_8_3_3;
  (* src = "crypto_accelerator.v:3319" *)
  input [7:0] io_keys_9_0_0;
  (* src = "crypto_accelerator.v:3320" *)
  input [7:0] io_keys_9_0_1;
  (* src = "crypto_accelerator.v:3321" *)
  input [7:0] io_keys_9_0_2;
  (* src = "crypto_accelerator.v:3322" *)
  input [7:0] io_keys_9_0_3;
  (* src = "crypto_accelerator.v:3323" *)
  input [7:0] io_keys_9_1_0;
  (* src = "crypto_accelerator.v:3324" *)
  input [7:0] io_keys_9_1_1;
  (* src = "crypto_accelerator.v:3325" *)
  input [7:0] io_keys_9_1_2;
  (* src = "crypto_accelerator.v:3326" *)
  input [7:0] io_keys_9_1_3;
  (* src = "crypto_accelerator.v:3327" *)
  input [7:0] io_keys_9_2_0;
  (* src = "crypto_accelerator.v:3328" *)
  input [7:0] io_keys_9_2_1;
  (* src = "crypto_accelerator.v:3329" *)
  input [7:0] io_keys_9_2_2;
  (* src = "crypto_accelerator.v:3330" *)
  input [7:0] io_keys_9_2_3;
  (* src = "crypto_accelerator.v:3331" *)
  input [7:0] io_keys_9_3_0;
  (* src = "crypto_accelerator.v:3332" *)
  input [7:0] io_keys_9_3_1;
  (* src = "crypto_accelerator.v:3333" *)
  input [7:0] io_keys_9_3_2;
  (* src = "crypto_accelerator.v:3334" *)
  input [7:0] io_keys_9_3_3;
  (* src = "crypto_accelerator.v:3422" *)
  output io_outputValid;
  (* src = "crypto_accelerator.v:3419" *)
  output io_ready;
  (* src = "crypto_accelerator.v:3418" *)
  output io_shift;
  (* src = "crypto_accelerator.v:3416" *)
  output io_shiftCyc;
  (* src = "crypto_accelerator.v:3417" *)
  output io_shiftRev;
  wire [2:0] keyEndAddr;
  (* src = "crypto_accelerator.v:3480" *)
  reg [7:0] matrix_0_0;
  (* src = "crypto_accelerator.v:3481" *)
  reg [7:0] matrix_0_1;
  (* src = "crypto_accelerator.v:3482" *)
  reg [7:0] matrix_0_2;
  (* src = "crypto_accelerator.v:3483" *)
  reg [7:0] matrix_0_3;
  (* src = "crypto_accelerator.v:3484" *)
  reg [7:0] matrix_1_0;
  (* src = "crypto_accelerator.v:3485" *)
  reg [7:0] matrix_1_1;
  (* src = "crypto_accelerator.v:3486" *)
  reg [7:0] matrix_1_2;
  (* src = "crypto_accelerator.v:3487" *)
  reg [7:0] matrix_1_3;
  (* src = "crypto_accelerator.v:3488" *)
  reg [7:0] matrix_2_0;
  (* src = "crypto_accelerator.v:3489" *)
  reg [7:0] matrix_2_1;
  (* src = "crypto_accelerator.v:3490" *)
  reg [7:0] matrix_2_2;
  (* src = "crypto_accelerator.v:3491" *)
  reg [7:0] matrix_2_3;
  (* src = "crypto_accelerator.v:3492" *)
  reg [7:0] matrix_3_0;
  (* src = "crypto_accelerator.v:3493" *)
  reg [7:0] matrix_3_1;
  (* src = "crypto_accelerator.v:3494" *)
  reg [7:0] matrix_3_2;
  (* src = "crypto_accelerator.v:3495" *)
  reg [7:0] matrix_3_3;
  (* src = "crypto_accelerator.v:3171" *)
  input reset;
  (* src = "crypto_accelerator.v:3635" *)
  wire [7:0] roundPart1_0_0;
  (* src = "crypto_accelerator.v:3773" *)
  wire [7:0] roundPart1_0_1;
  (* src = "crypto_accelerator.v:3911" *)
  wire [7:0] roundPart1_0_2;
  (* src = "crypto_accelerator.v:4049" *)
  wire [7:0] roundPart1_0_3;
  (* src = "crypto_accelerator.v:4187" *)
  wire [7:0] roundPart1_1_0;
  (* src = "crypto_accelerator.v:4325" *)
  wire [7:0] roundPart1_1_1;
  (* src = "crypto_accelerator.v:4463" *)
  wire [7:0] roundPart1_1_2;
  (* src = "crypto_accelerator.v:4601" *)
  wire [7:0] roundPart1_1_3;
  (* src = "crypto_accelerator.v:4739" *)
  wire [7:0] roundPart1_2_0;
  (* src = "crypto_accelerator.v:4877" *)
  wire [7:0] roundPart1_2_1;
  (* src = "crypto_accelerator.v:5015" *)
  wire [7:0] roundPart1_2_2;
  (* src = "crypto_accelerator.v:5153" *)
  wire [7:0] roundPart1_2_3;
  (* src = "crypto_accelerator.v:5291" *)
  wire [7:0] roundPart1_3_0;
  (* src = "crypto_accelerator.v:5429" *)
  wire [7:0] roundPart1_3_1;
  (* src = "crypto_accelerator.v:5567" *)
  wire [7:0] roundPart1_3_2;
  (* src = "crypto_accelerator.v:5705" *)
  wire [7:0] roundPart1_3_3;
  (* src = "crypto_accelerator.v:3476" *)
  reg [5:0] state;
  (* src = "crypto_accelerator.v:5931" *)
  wire [7:0] xorOut_0_0;
  (* src = "crypto_accelerator.v:5932" *)
  wire [7:0] xorOut_0_1;
  (* src = "crypto_accelerator.v:5933" *)
  wire [7:0] xorOut_0_2;
  (* src = "crypto_accelerator.v:5934" *)
  wire [7:0] xorOut_0_3;
  (* src = "crypto_accelerator.v:5935" *)
  wire [7:0] xorOut_1_0;
  (* src = "crypto_accelerator.v:5936" *)
  wire [7:0] xorOut_1_1;
  (* src = "crypto_accelerator.v:5937" *)
  wire [7:0] xorOut_1_2;
  (* src = "crypto_accelerator.v:5938" *)
  wire [7:0] xorOut_1_3;
  (* src = "crypto_accelerator.v:5939" *)
  wire [7:0] xorOut_2_0;
  (* src = "crypto_accelerator.v:5940" *)
  wire [7:0] xorOut_2_1;
  (* src = "crypto_accelerator.v:5941" *)
  wire [7:0] xorOut_2_2;
  (* src = "crypto_accelerator.v:5942" *)
  wire [7:0] xorOut_2_3;
  (* src = "crypto_accelerator.v:5943" *)
  wire [7:0] xorOut_3_0;
  (* src = "crypto_accelerator.v:5944" *)
  wire [7:0] xorOut_3_1;
  (* src = "crypto_accelerator.v:5945" *)
  wire [7:0] xorOut_3_2;
  (* src = "crypto_accelerator.v:5946" *)
  wire [7:0] xorOut_3_3;
  assign _T_105 = _T_66 & (* src = "crypto_accelerator.v:3535" *) _T_93;
  assign _T_107 = _T_41 & (* src = "crypto_accelerator.v:3536" *) _T_57;
  assign _T_111 = _T_59 & (* src = "crypto_accelerator.v:3538" *) _T_91;
  assign _T_115 = _T_68 & (* src = "crypto_accelerator.v:3540" *) _T_95;
  assign _T_117 = _T_44 & (* src = "crypto_accelerator.v:3541" *) _T_62;
  assign _T_121 = _T_78 & (* src = "crypto_accelerator.v:3543" *) _T_76;
  assign _T_125 = _T_49 & (* src = "crypto_accelerator.v:3545" *) _T_99;
  assign _T_127 = _T_80 & (* src = "crypto_accelerator.v:3546" *) _T_97;
  assign _T_131 = _T_47 & (* src = "crypto_accelerator.v:3548" *) _T_64;
  assign _T_153 = _T_147 & (* src = "crypto_accelerator.v:3559" *) _T_143;
  assign _T_161 = _T_159 & (* src = "crypto_accelerator.v:3563" *) _T_157;
  assign _T_163 = _T_155 & (* src = "crypto_accelerator.v:3564" *) _T_151;
  assign _T_165 = _T_143 & (* src = "crypto_accelerator.v:3565" *) _T_149;
  assign _T_167 = _T_157 & (* src = "crypto_accelerator.v:3566" *) _T_165;
  assign _T_171 = _T_145 & (* src = "crypto_accelerator.v:3568" *) _T_147;
  assign _T_173 = _T_151 & (* src = "crypto_accelerator.v:3569" *) _T_171;
  assign _T_195 = _T_191 & (* src = "crypto_accelerator.v:3580" *) _T_93;
  assign _T_197 = _T_183 & (* src = "crypto_accelerator.v:3581" *) _T_57;
  assign _T_199 = _T_181 & (* src = "crypto_accelerator.v:3582" *) _T_91;
  assign _T_201 = _T_189 & (* src = "crypto_accelerator.v:3583" *) _T_95;
  assign _T_203 = _T_179 & (* src = "crypto_accelerator.v:3584" *) _T_62;
  assign _T_205 = _T_177 & (* src = "crypto_accelerator.v:3585" *) _T_76;
  assign _T_207 = _T_187 & (* src = "crypto_accelerator.v:3586" *) _T_99;
  assign _T_209 = _T_193 & (* src = "crypto_accelerator.v:3587" *) _T_97;
  assign _T_211 = _T_185 & (* src = "crypto_accelerator.v:3588" *) _T_64;
  assign _T_213 = _T_191 & (* src = "crypto_accelerator.v:3589" *) _T_66;
  assign _T_215 = _T_183 & (* src = "crypto_accelerator.v:3590" *) _T_41;
  assign _T_217 = _T_181 & (* src = "crypto_accelerator.v:3591" *) _T_59;
  assign _T_219 = _T_189 & (* src = "crypto_accelerator.v:3592" *) _T_68;
  assign _T_221 = _T_179 & (* src = "crypto_accelerator.v:3593" *) _T_44;
  assign _T_223 = _T_177 & (* src = "crypto_accelerator.v:3594" *) _T_78;
  assign _T_225 = _T_187 & (* src = "crypto_accelerator.v:3595" *) _T_49;
  assign _T_227 = _T_193 & (* src = "crypto_accelerator.v:3596" *) _T_80;
  assign _T_229 = _T_185 & (* src = "crypto_accelerator.v:3597" *) _T_47;
  assign _T_384 = _T_345 & (* src = "crypto_accelerator.v:3673" *) _T_372;
  assign _T_386 = _T_320 & (* src = "crypto_accelerator.v:3674" *) _T_336;
  assign _T_390 = _T_338 & (* src = "crypto_accelerator.v:3676" *) _T_370;
  assign _T_394 = _T_347 & (* src = "crypto_accelerator.v:3678" *) _T_374;
  assign _T_396 = _T_323 & (* src = "crypto_accelerator.v:3679" *) _T_341;
  assign _T_400 = _T_357 & (* src = "crypto_accelerator.v:3681" *) _T_355;
  assign _T_404 = _T_328 & (* src = "crypto_accelerator.v:3683" *) _T_378;
  assign _T_406 = _T_359 & (* src = "crypto_accelerator.v:3684" *) _T_376;
  assign _T_410 = _T_326 & (* src = "crypto_accelerator.v:3686" *) _T_343;
  assign _T_432 = _T_426 & (* src = "crypto_accelerator.v:3697" *) _T_422;
  assign _T_440 = _T_438 & (* src = "crypto_accelerator.v:3701" *) _T_436;
  assign _T_442 = _T_434 & (* src = "crypto_accelerator.v:3702" *) _T_430;
  assign _T_444 = _T_422 & (* src = "crypto_accelerator.v:3703" *) _T_428;
  assign _T_446 = _T_436 & (* src = "crypto_accelerator.v:3704" *) _T_444;
  assign _T_450 = _T_424 & (* src = "crypto_accelerator.v:3706" *) _T_426;
  assign _T_452 = _T_430 & (* src = "crypto_accelerator.v:3707" *) _T_450;
  assign _T_474 = _T_470 & (* src = "crypto_accelerator.v:3718" *) _T_372;
  assign _T_476 = _T_462 & (* src = "crypto_accelerator.v:3719" *) _T_336;
  assign _T_478 = _T_460 & (* src = "crypto_accelerator.v:3720" *) _T_370;
  assign _T_480 = _T_468 & (* src = "crypto_accelerator.v:3721" *) _T_374;
  assign _T_482 = _T_458 & (* src = "crypto_accelerator.v:3722" *) _T_341;
  assign _T_484 = _T_456 & (* src = "crypto_accelerator.v:3723" *) _T_355;
  assign _T_486 = _T_466 & (* src = "crypto_accelerator.v:3724" *) _T_378;
  assign _T_488 = _T_472 & (* src = "crypto_accelerator.v:3725" *) _T_376;
  assign _T_490 = _T_464 & (* src = "crypto_accelerator.v:3726" *) _T_343;
  assign _T_492 = _T_470 & (* src = "crypto_accelerator.v:3727" *) _T_345;
  assign _T_494 = _T_462 & (* src = "crypto_accelerator.v:3728" *) _T_320;
  assign _T_496 = _T_460 & (* src = "crypto_accelerator.v:3729" *) _T_338;
  assign _T_498 = _T_468 & (* src = "crypto_accelerator.v:3730" *) _T_347;
  assign _T_500 = _T_458 & (* src = "crypto_accelerator.v:3731" *) _T_323;
  assign _T_502 = _T_456 & (* src = "crypto_accelerator.v:3732" *) _T_357;
  assign _T_504 = _T_466 & (* src = "crypto_accelerator.v:3733" *) _T_328;
  assign _T_506 = _T_472 & (* src = "crypto_accelerator.v:3734" *) _T_359;
  assign _T_508 = _T_464 & (* src = "crypto_accelerator.v:3735" *) _T_326;
  assign _T_663 = _T_624 & (* src = "crypto_accelerator.v:3811" *) _T_651;
  assign _T_665 = _T_599 & (* src = "crypto_accelerator.v:3812" *) _T_615;
  assign _T_669 = _T_617 & (* src = "crypto_accelerator.v:3814" *) _T_649;
  assign _T_673 = _T_626 & (* src = "crypto_accelerator.v:3816" *) _T_653;
  assign _T_675 = _T_602 & (* src = "crypto_accelerator.v:3817" *) _T_620;
  assign _T_679 = _T_636 & (* src = "crypto_accelerator.v:3819" *) _T_634;
  assign _T_683 = _T_607 & (* src = "crypto_accelerator.v:3821" *) _T_657;
  assign _T_685 = _T_638 & (* src = "crypto_accelerator.v:3822" *) _T_655;
  assign _T_689 = _T_605 & (* src = "crypto_accelerator.v:3824" *) _T_622;
  assign _T_711 = _T_705 & (* src = "crypto_accelerator.v:3835" *) _T_701;
  assign _T_719 = _T_717 & (* src = "crypto_accelerator.v:3839" *) _T_715;
  assign _T_721 = _T_713 & (* src = "crypto_accelerator.v:3840" *) _T_709;
  assign _T_723 = _T_701 & (* src = "crypto_accelerator.v:3841" *) _T_707;
  assign _T_725 = _T_715 & (* src = "crypto_accelerator.v:3842" *) _T_723;
  assign _T_729 = _T_703 & (* src = "crypto_accelerator.v:3844" *) _T_705;
  assign _T_731 = _T_709 & (* src = "crypto_accelerator.v:3845" *) _T_729;
  assign _T_753 = _T_749 & (* src = "crypto_accelerator.v:3856" *) _T_651;
  assign _T_755 = _T_741 & (* src = "crypto_accelerator.v:3857" *) _T_615;
  assign _T_757 = _T_739 & (* src = "crypto_accelerator.v:3858" *) _T_649;
  assign _T_759 = _T_747 & (* src = "crypto_accelerator.v:3859" *) _T_653;
  assign _T_761 = _T_737 & (* src = "crypto_accelerator.v:3860" *) _T_620;
  assign _T_763 = _T_735 & (* src = "crypto_accelerator.v:3861" *) _T_634;
  assign _T_765 = _T_745 & (* src = "crypto_accelerator.v:3862" *) _T_657;
  assign _T_767 = _T_751 & (* src = "crypto_accelerator.v:3863" *) _T_655;
  assign _T_769 = _T_743 & (* src = "crypto_accelerator.v:3864" *) _T_622;
  assign _T_771 = _T_749 & (* src = "crypto_accelerator.v:3865" *) _T_624;
  assign _T_773 = _T_741 & (* src = "crypto_accelerator.v:3866" *) _T_599;
  assign _T_775 = _T_739 & (* src = "crypto_accelerator.v:3867" *) _T_617;
  assign _T_777 = _T_747 & (* src = "crypto_accelerator.v:3868" *) _T_626;
  assign _T_779 = _T_737 & (* src = "crypto_accelerator.v:3869" *) _T_602;
  assign _T_781 = _T_735 & (* src = "crypto_accelerator.v:3870" *) _T_636;
  assign _T_783 = _T_745 & (* src = "crypto_accelerator.v:3871" *) _T_607;
  assign _T_785 = _T_751 & (* src = "crypto_accelerator.v:3872" *) _T_638;
  assign _T_787 = _T_743 & (* src = "crypto_accelerator.v:3873" *) _T_605;
  assign _T_942 = _T_903 & (* src = "crypto_accelerator.v:3949" *) _T_930;
  assign _T_944 = _T_878 & (* src = "crypto_accelerator.v:3950" *) _T_894;
  assign _T_948 = _T_896 & (* src = "crypto_accelerator.v:3952" *) _T_928;
  assign _T_952 = _T_905 & (* src = "crypto_accelerator.v:3954" *) _T_932;
  assign _T_954 = _T_881 & (* src = "crypto_accelerator.v:3955" *) _T_899;
  assign _T_958 = _T_915 & (* src = "crypto_accelerator.v:3957" *) _T_913;
  assign _T_962 = _T_886 & (* src = "crypto_accelerator.v:3959" *) _T_936;
  assign _T_964 = _T_917 & (* src = "crypto_accelerator.v:3960" *) _T_934;
  assign _T_968 = _T_884 & (* src = "crypto_accelerator.v:3962" *) _T_901;
  assign _T_990 = _T_984 & (* src = "crypto_accelerator.v:3973" *) _T_980;
  assign _T_998 = _T_996 & (* src = "crypto_accelerator.v:3977" *) _T_994;
  assign _T_1000 = _T_992 & (* src = "crypto_accelerator.v:3978" *) _T_988;
  assign _T_1002 = _T_980 & (* src = "crypto_accelerator.v:3979" *) _T_986;
  assign _T_1004 = _T_994 & (* src = "crypto_accelerator.v:3980" *) _T_1002;
  assign _T_1008 = _T_982 & (* src = "crypto_accelerator.v:3982" *) _T_984;
  assign _T_1010 = _T_988 & (* src = "crypto_accelerator.v:3983" *) _T_1008;
  assign _T_1032 = _T_1028 & (* src = "crypto_accelerator.v:3994" *) _T_930;
  assign _T_1034 = _T_1020 & (* src = "crypto_accelerator.v:3995" *) _T_894;
  assign _T_1036 = _T_1018 & (* src = "crypto_accelerator.v:3996" *) _T_928;
  assign _T_1038 = _T_1026 & (* src = "crypto_accelerator.v:3997" *) _T_932;
  assign _T_1040 = _T_1016 & (* src = "crypto_accelerator.v:3998" *) _T_899;
  assign _T_1042 = _T_1014 & (* src = "crypto_accelerator.v:3999" *) _T_913;
  assign _T_1044 = _T_1024 & (* src = "crypto_accelerator.v:4000" *) _T_936;
  assign _T_1046 = _T_1030 & (* src = "crypto_accelerator.v:4001" *) _T_934;
  assign _T_1048 = _T_1022 & (* src = "crypto_accelerator.v:4002" *) _T_901;
  assign _T_1050 = _T_1028 & (* src = "crypto_accelerator.v:4003" *) _T_903;
  assign _T_1052 = _T_1020 & (* src = "crypto_accelerator.v:4004" *) _T_878;
  assign _T_1054 = _T_1018 & (* src = "crypto_accelerator.v:4005" *) _T_896;
  assign _T_1056 = _T_1026 & (* src = "crypto_accelerator.v:4006" *) _T_905;
  assign _T_1058 = _T_1016 & (* src = "crypto_accelerator.v:4007" *) _T_881;
  assign _T_1060 = _T_1014 & (* src = "crypto_accelerator.v:4008" *) _T_915;
  assign _T_1062 = _T_1024 & (* src = "crypto_accelerator.v:4009" *) _T_886;
  assign _T_1064 = _T_1030 & (* src = "crypto_accelerator.v:4010" *) _T_917;
  assign _T_1066 = _T_1022 & (* src = "crypto_accelerator.v:4011" *) _T_884;
  assign _T_1222 = _T_1183 & (* src = "crypto_accelerator.v:4087" *) _T_1210;
  assign _T_1224 = _T_1158 & (* src = "crypto_accelerator.v:4088" *) _T_1174;
  assign _T_1228 = _T_1176 & (* src = "crypto_accelerator.v:4090" *) _T_1208;
  assign _T_1232 = _T_1185 & (* src = "crypto_accelerator.v:4092" *) _T_1212;
  assign _T_1234 = _T_1161 & (* src = "crypto_accelerator.v:4093" *) _T_1179;
  assign _T_1238 = _T_1195 & (* src = "crypto_accelerator.v:4095" *) _T_1193;
  assign _T_1242 = _T_1166 & (* src = "crypto_accelerator.v:4097" *) _T_1216;
  assign _T_1244 = _T_1197 & (* src = "crypto_accelerator.v:4098" *) _T_1214;
  assign _T_1248 = _T_1164 & (* src = "crypto_accelerator.v:4100" *) _T_1181;
  assign _T_1270 = _T_1264 & (* src = "crypto_accelerator.v:4111" *) _T_1260;
  assign _T_1278 = _T_1276 & (* src = "crypto_accelerator.v:4115" *) _T_1274;
  assign _T_1280 = _T_1272 & (* src = "crypto_accelerator.v:4116" *) _T_1268;
  assign _T_1282 = _T_1260 & (* src = "crypto_accelerator.v:4117" *) _T_1266;
  assign _T_1284 = _T_1274 & (* src = "crypto_accelerator.v:4118" *) _T_1282;
  assign _T_1288 = _T_1262 & (* src = "crypto_accelerator.v:4120" *) _T_1264;
  assign _T_1290 = _T_1268 & (* src = "crypto_accelerator.v:4121" *) _T_1288;
  assign _T_1312 = _T_1308 & (* src = "crypto_accelerator.v:4132" *) _T_1210;
  assign _T_1314 = _T_1300 & (* src = "crypto_accelerator.v:4133" *) _T_1174;
  assign _T_1316 = _T_1298 & (* src = "crypto_accelerator.v:4134" *) _T_1208;
  assign _T_1318 = _T_1306 & (* src = "crypto_accelerator.v:4135" *) _T_1212;
  assign _T_1320 = _T_1296 & (* src = "crypto_accelerator.v:4136" *) _T_1179;
  assign _T_1322 = _T_1294 & (* src = "crypto_accelerator.v:4137" *) _T_1193;
  assign _T_1324 = _T_1304 & (* src = "crypto_accelerator.v:4138" *) _T_1216;
  assign _T_1326 = _T_1310 & (* src = "crypto_accelerator.v:4139" *) _T_1214;
  assign _T_1328 = _T_1302 & (* src = "crypto_accelerator.v:4140" *) _T_1181;
  assign _T_1330 = _T_1308 & (* src = "crypto_accelerator.v:4141" *) _T_1183;
  assign _T_1332 = _T_1300 & (* src = "crypto_accelerator.v:4142" *) _T_1158;
  assign _T_1334 = _T_1298 & (* src = "crypto_accelerator.v:4143" *) _T_1176;
  assign _T_1336 = _T_1306 & (* src = "crypto_accelerator.v:4144" *) _T_1185;
  assign _T_1338 = _T_1296 & (* src = "crypto_accelerator.v:4145" *) _T_1161;
  assign _T_1340 = _T_1294 & (* src = "crypto_accelerator.v:4146" *) _T_1195;
  assign _T_1342 = _T_1304 & (* src = "crypto_accelerator.v:4147" *) _T_1166;
  assign _T_1344 = _T_1310 & (* src = "crypto_accelerator.v:4148" *) _T_1197;
  assign _T_1346 = _T_1302 & (* src = "crypto_accelerator.v:4149" *) _T_1164;
  assign _T_1501 = _T_1462 & (* src = "crypto_accelerator.v:4225" *) _T_1489;
  assign _T_1503 = _T_1437 & (* src = "crypto_accelerator.v:4226" *) _T_1453;
  assign _T_1507 = _T_1455 & (* src = "crypto_accelerator.v:4228" *) _T_1487;
  assign _T_1511 = _T_1464 & (* src = "crypto_accelerator.v:4230" *) _T_1491;
  assign _T_1513 = _T_1440 & (* src = "crypto_accelerator.v:4231" *) _T_1458;
  assign _T_1517 = _T_1474 & (* src = "crypto_accelerator.v:4233" *) _T_1472;
  assign _T_1521 = _T_1445 & (* src = "crypto_accelerator.v:4235" *) _T_1495;
  assign _T_1523 = _T_1476 & (* src = "crypto_accelerator.v:4236" *) _T_1493;
  assign _T_1527 = _T_1443 & (* src = "crypto_accelerator.v:4238" *) _T_1460;
  assign _T_1549 = _T_1543 & (* src = "crypto_accelerator.v:4249" *) _T_1539;
  assign _T_1557 = _T_1555 & (* src = "crypto_accelerator.v:4253" *) _T_1553;
  assign _T_1559 = _T_1551 & (* src = "crypto_accelerator.v:4254" *) _T_1547;
  assign _T_1561 = _T_1539 & (* src = "crypto_accelerator.v:4255" *) _T_1545;
  assign _T_1563 = _T_1553 & (* src = "crypto_accelerator.v:4256" *) _T_1561;
  assign _T_1567 = _T_1541 & (* src = "crypto_accelerator.v:4258" *) _T_1543;
  assign _T_1569 = _T_1547 & (* src = "crypto_accelerator.v:4259" *) _T_1567;
  assign _T_1591 = _T_1587 & (* src = "crypto_accelerator.v:4270" *) _T_1489;
  assign _T_1593 = _T_1579 & (* src = "crypto_accelerator.v:4271" *) _T_1453;
  assign _T_1595 = _T_1577 & (* src = "crypto_accelerator.v:4272" *) _T_1487;
  assign _T_1597 = _T_1585 & (* src = "crypto_accelerator.v:4273" *) _T_1491;
  assign _T_1599 = _T_1575 & (* src = "crypto_accelerator.v:4274" *) _T_1458;
  assign _T_1601 = _T_1573 & (* src = "crypto_accelerator.v:4275" *) _T_1472;
  assign _T_1603 = _T_1583 & (* src = "crypto_accelerator.v:4276" *) _T_1495;
  assign _T_1605 = _T_1589 & (* src = "crypto_accelerator.v:4277" *) _T_1493;
  assign _T_1607 = _T_1581 & (* src = "crypto_accelerator.v:4278" *) _T_1460;
  assign _T_1609 = _T_1587 & (* src = "crypto_accelerator.v:4279" *) _T_1462;
  assign _T_1611 = _T_1579 & (* src = "crypto_accelerator.v:4280" *) _T_1437;
  assign _T_1613 = _T_1577 & (* src = "crypto_accelerator.v:4281" *) _T_1455;
  assign _T_1615 = _T_1585 & (* src = "crypto_accelerator.v:4282" *) _T_1464;
  assign _T_1617 = _T_1575 & (* src = "crypto_accelerator.v:4283" *) _T_1440;
  assign _T_1619 = _T_1573 & (* src = "crypto_accelerator.v:4284" *) _T_1474;
  assign _T_1621 = _T_1583 & (* src = "crypto_accelerator.v:4285" *) _T_1445;
  assign _T_1623 = _T_1589 & (* src = "crypto_accelerator.v:4286" *) _T_1476;
  assign _T_1625 = _T_1581 & (* src = "crypto_accelerator.v:4287" *) _T_1443;
  assign _T_1780 = _T_1741 & (* src = "crypto_accelerator.v:4363" *) _T_1768;
  assign _T_1782 = _T_1716 & (* src = "crypto_accelerator.v:4364" *) _T_1732;
  assign _T_1786 = _T_1734 & (* src = "crypto_accelerator.v:4366" *) _T_1766;
  assign _T_1790 = _T_1743 & (* src = "crypto_accelerator.v:4368" *) _T_1770;
  assign _T_1792 = _T_1719 & (* src = "crypto_accelerator.v:4369" *) _T_1737;
  assign _T_1796 = _T_1753 & (* src = "crypto_accelerator.v:4371" *) _T_1751;
  assign _T_1800 = _T_1724 & (* src = "crypto_accelerator.v:4373" *) _T_1774;
  assign _T_1802 = _T_1755 & (* src = "crypto_accelerator.v:4374" *) _T_1772;
  assign _T_1806 = _T_1722 & (* src = "crypto_accelerator.v:4376" *) _T_1739;
  assign _T_1828 = _T_1822 & (* src = "crypto_accelerator.v:4387" *) _T_1818;
  assign _T_1836 = _T_1834 & (* src = "crypto_accelerator.v:4391" *) _T_1832;
  assign _T_1838 = _T_1830 & (* src = "crypto_accelerator.v:4392" *) _T_1826;
  assign _T_1840 = _T_1818 & (* src = "crypto_accelerator.v:4393" *) _T_1824;
  assign _T_1842 = _T_1832 & (* src = "crypto_accelerator.v:4394" *) _T_1840;
  assign _T_1846 = _T_1820 & (* src = "crypto_accelerator.v:4396" *) _T_1822;
  assign _T_1848 = _T_1826 & (* src = "crypto_accelerator.v:4397" *) _T_1846;
  assign _T_1870 = _T_1866 & (* src = "crypto_accelerator.v:4408" *) _T_1768;
  assign _T_1872 = _T_1858 & (* src = "crypto_accelerator.v:4409" *) _T_1732;
  assign _T_1874 = _T_1856 & (* src = "crypto_accelerator.v:4410" *) _T_1766;
  assign _T_1876 = _T_1864 & (* src = "crypto_accelerator.v:4411" *) _T_1770;
  assign _T_1878 = _T_1854 & (* src = "crypto_accelerator.v:4412" *) _T_1737;
  assign _T_1880 = _T_1852 & (* src = "crypto_accelerator.v:4413" *) _T_1751;
  assign _T_1882 = _T_1862 & (* src = "crypto_accelerator.v:4414" *) _T_1774;
  assign _T_1884 = _T_1868 & (* src = "crypto_accelerator.v:4415" *) _T_1772;
  assign _T_1886 = _T_1860 & (* src = "crypto_accelerator.v:4416" *) _T_1739;
  assign _T_1888 = _T_1866 & (* src = "crypto_accelerator.v:4417" *) _T_1741;
  assign _T_1890 = _T_1858 & (* src = "crypto_accelerator.v:4418" *) _T_1716;
  assign _T_1892 = _T_1856 & (* src = "crypto_accelerator.v:4419" *) _T_1734;
  assign _T_1894 = _T_1864 & (* src = "crypto_accelerator.v:4420" *) _T_1743;
  assign _T_1896 = _T_1854 & (* src = "crypto_accelerator.v:4421" *) _T_1719;
  assign _T_1898 = _T_1852 & (* src = "crypto_accelerator.v:4422" *) _T_1753;
  assign _T_1900 = _T_1862 & (* src = "crypto_accelerator.v:4423" *) _T_1724;
  assign _T_1902 = _T_1868 & (* src = "crypto_accelerator.v:4424" *) _T_1755;
  assign _T_1904 = _T_1860 & (* src = "crypto_accelerator.v:4425" *) _T_1722;
  assign _T_2059 = _T_2020 & (* src = "crypto_accelerator.v:4501" *) _T_2047;
  assign _T_2061 = _T_1995 & (* src = "crypto_accelerator.v:4502" *) _T_2011;
  assign _T_2065 = _T_2013 & (* src = "crypto_accelerator.v:4504" *) _T_2045;
  assign _T_2069 = _T_2022 & (* src = "crypto_accelerator.v:4506" *) _T_2049;
  assign _T_2071 = _T_1998 & (* src = "crypto_accelerator.v:4507" *) _T_2016;
  assign _T_2075 = _T_2032 & (* src = "crypto_accelerator.v:4509" *) _T_2030;
  assign _T_2079 = _T_2003 & (* src = "crypto_accelerator.v:4511" *) _T_2053;
  assign _T_2081 = _T_2034 & (* src = "crypto_accelerator.v:4512" *) _T_2051;
  assign _T_2085 = _T_2001 & (* src = "crypto_accelerator.v:4514" *) _T_2018;
  assign _T_2107 = _T_2101 & (* src = "crypto_accelerator.v:4525" *) _T_2097;
  assign _T_2115 = _T_2113 & (* src = "crypto_accelerator.v:4529" *) _T_2111;
  assign _T_2117 = _T_2109 & (* src = "crypto_accelerator.v:4530" *) _T_2105;
  assign _T_2119 = _T_2097 & (* src = "crypto_accelerator.v:4531" *) _T_2103;
  assign _T_2121 = _T_2111 & (* src = "crypto_accelerator.v:4532" *) _T_2119;
  assign _T_2125 = _T_2099 & (* src = "crypto_accelerator.v:4534" *) _T_2101;
  assign _T_2127 = _T_2105 & (* src = "crypto_accelerator.v:4535" *) _T_2125;
  assign _T_2149 = _T_2145 & (* src = "crypto_accelerator.v:4546" *) _T_2047;
  assign _T_2151 = _T_2137 & (* src = "crypto_accelerator.v:4547" *) _T_2011;
  assign _T_2153 = _T_2135 & (* src = "crypto_accelerator.v:4548" *) _T_2045;
  assign _T_2155 = _T_2143 & (* src = "crypto_accelerator.v:4549" *) _T_2049;
  assign _T_2157 = _T_2133 & (* src = "crypto_accelerator.v:4550" *) _T_2016;
  assign _T_2159 = _T_2131 & (* src = "crypto_accelerator.v:4551" *) _T_2030;
  assign _T_2161 = _T_2141 & (* src = "crypto_accelerator.v:4552" *) _T_2053;
  assign _T_2163 = _T_2147 & (* src = "crypto_accelerator.v:4553" *) _T_2051;
  assign _T_2165 = _T_2139 & (* src = "crypto_accelerator.v:4554" *) _T_2018;
  assign _T_2167 = _T_2145 & (* src = "crypto_accelerator.v:4555" *) _T_2020;
  assign _T_2169 = _T_2137 & (* src = "crypto_accelerator.v:4556" *) _T_1995;
  assign _T_2171 = _T_2135 & (* src = "crypto_accelerator.v:4557" *) _T_2013;
  assign _T_2173 = _T_2143 & (* src = "crypto_accelerator.v:4558" *) _T_2022;
  assign _T_2175 = _T_2133 & (* src = "crypto_accelerator.v:4559" *) _T_1998;
  assign _T_2177 = _T_2131 & (* src = "crypto_accelerator.v:4560" *) _T_2032;
  assign _T_2179 = _T_2141 & (* src = "crypto_accelerator.v:4561" *) _T_2003;
  assign _T_2181 = _T_2147 & (* src = "crypto_accelerator.v:4562" *) _T_2034;
  assign _T_2183 = _T_2139 & (* src = "crypto_accelerator.v:4563" *) _T_2001;
  assign _T_2339 = _T_2300 & (* src = "crypto_accelerator.v:4639" *) _T_2327;
  assign _T_2341 = _T_2275 & (* src = "crypto_accelerator.v:4640" *) _T_2291;
  assign _T_2345 = _T_2293 & (* src = "crypto_accelerator.v:4642" *) _T_2325;
  assign _T_2349 = _T_2302 & (* src = "crypto_accelerator.v:4644" *) _T_2329;
  assign _T_2351 = _T_2278 & (* src = "crypto_accelerator.v:4645" *) _T_2296;
  assign _T_2355 = _T_2312 & (* src = "crypto_accelerator.v:4647" *) _T_2310;
  assign _T_2359 = _T_2283 & (* src = "crypto_accelerator.v:4649" *) _T_2333;
  assign _T_2361 = _T_2314 & (* src = "crypto_accelerator.v:4650" *) _T_2331;
  assign _T_2365 = _T_2281 & (* src = "crypto_accelerator.v:4652" *) _T_2298;
  assign _T_2387 = _T_2381 & (* src = "crypto_accelerator.v:4663" *) _T_2377;
  assign _T_2395 = _T_2393 & (* src = "crypto_accelerator.v:4667" *) _T_2391;
  assign _T_2397 = _T_2389 & (* src = "crypto_accelerator.v:4668" *) _T_2385;
  assign _T_2399 = _T_2377 & (* src = "crypto_accelerator.v:4669" *) _T_2383;
  assign _T_2401 = _T_2391 & (* src = "crypto_accelerator.v:4670" *) _T_2399;
  assign _T_2405 = _T_2379 & (* src = "crypto_accelerator.v:4672" *) _T_2381;
  assign _T_2407 = _T_2385 & (* src = "crypto_accelerator.v:4673" *) _T_2405;
  assign _T_2429 = _T_2425 & (* src = "crypto_accelerator.v:4684" *) _T_2327;
  assign _T_2431 = _T_2417 & (* src = "crypto_accelerator.v:4685" *) _T_2291;
  assign _T_2433 = _T_2415 & (* src = "crypto_accelerator.v:4686" *) _T_2325;
  assign _T_2435 = _T_2423 & (* src = "crypto_accelerator.v:4687" *) _T_2329;
  assign _T_2437 = _T_2413 & (* src = "crypto_accelerator.v:4688" *) _T_2296;
  assign _T_2439 = _T_2411 & (* src = "crypto_accelerator.v:4689" *) _T_2310;
  assign _T_2441 = _T_2421 & (* src = "crypto_accelerator.v:4690" *) _T_2333;
  assign _T_2443 = _T_2427 & (* src = "crypto_accelerator.v:4691" *) _T_2331;
  assign _T_2445 = _T_2419 & (* src = "crypto_accelerator.v:4692" *) _T_2298;
  assign _T_2447 = _T_2425 & (* src = "crypto_accelerator.v:4693" *) _T_2300;
  assign _T_2449 = _T_2417 & (* src = "crypto_accelerator.v:4694" *) _T_2275;
  assign _T_2451 = _T_2415 & (* src = "crypto_accelerator.v:4695" *) _T_2293;
  assign _T_2453 = _T_2423 & (* src = "crypto_accelerator.v:4696" *) _T_2302;
  assign _T_2455 = _T_2413 & (* src = "crypto_accelerator.v:4697" *) _T_2278;
  assign _T_2457 = _T_2411 & (* src = "crypto_accelerator.v:4698" *) _T_2312;
  assign _T_2459 = _T_2421 & (* src = "crypto_accelerator.v:4699" *) _T_2283;
  assign _T_2461 = _T_2427 & (* src = "crypto_accelerator.v:4700" *) _T_2314;
  assign _T_2463 = _T_2419 & (* src = "crypto_accelerator.v:4701" *) _T_2281;
  assign _T_2618 = _T_2579 & (* src = "crypto_accelerator.v:4777" *) _T_2606;
  assign _T_2620 = _T_2554 & (* src = "crypto_accelerator.v:4778" *) _T_2570;
  assign _T_2624 = _T_2572 & (* src = "crypto_accelerator.v:4780" *) _T_2604;
  assign _T_2628 = _T_2581 & (* src = "crypto_accelerator.v:4782" *) _T_2608;
  assign _T_2630 = _T_2557 & (* src = "crypto_accelerator.v:4783" *) _T_2575;
  assign _T_2634 = _T_2591 & (* src = "crypto_accelerator.v:4785" *) _T_2589;
  assign _T_2638 = _T_2562 & (* src = "crypto_accelerator.v:4787" *) _T_2612;
  assign _T_2640 = _T_2593 & (* src = "crypto_accelerator.v:4788" *) _T_2610;
  assign _T_2644 = _T_2560 & (* src = "crypto_accelerator.v:4790" *) _T_2577;
  assign _T_2666 = _T_2660 & (* src = "crypto_accelerator.v:4801" *) _T_2656;
  assign _T_2674 = _T_2672 & (* src = "crypto_accelerator.v:4805" *) _T_2670;
  assign _T_2676 = _T_2668 & (* src = "crypto_accelerator.v:4806" *) _T_2664;
  assign _T_2678 = _T_2656 & (* src = "crypto_accelerator.v:4807" *) _T_2662;
  assign _T_2680 = _T_2670 & (* src = "crypto_accelerator.v:4808" *) _T_2678;
  assign _T_2684 = _T_2658 & (* src = "crypto_accelerator.v:4810" *) _T_2660;
  assign _T_2686 = _T_2664 & (* src = "crypto_accelerator.v:4811" *) _T_2684;
  assign _T_2708 = _T_2704 & (* src = "crypto_accelerator.v:4822" *) _T_2606;
  assign _T_2710 = _T_2696 & (* src = "crypto_accelerator.v:4823" *) _T_2570;
  assign _T_2712 = _T_2694 & (* src = "crypto_accelerator.v:4824" *) _T_2604;
  assign _T_2714 = _T_2702 & (* src = "crypto_accelerator.v:4825" *) _T_2608;
  assign _T_2716 = _T_2692 & (* src = "crypto_accelerator.v:4826" *) _T_2575;
  assign _T_2718 = _T_2690 & (* src = "crypto_accelerator.v:4827" *) _T_2589;
  assign _T_2720 = _T_2700 & (* src = "crypto_accelerator.v:4828" *) _T_2612;
  assign _T_2722 = _T_2706 & (* src = "crypto_accelerator.v:4829" *) _T_2610;
  assign _T_2724 = _T_2698 & (* src = "crypto_accelerator.v:4830" *) _T_2577;
  assign _T_2726 = _T_2704 & (* src = "crypto_accelerator.v:4831" *) _T_2579;
  assign _T_2728 = _T_2696 & (* src = "crypto_accelerator.v:4832" *) _T_2554;
  assign _T_2730 = _T_2694 & (* src = "crypto_accelerator.v:4833" *) _T_2572;
  assign _T_2732 = _T_2702 & (* src = "crypto_accelerator.v:4834" *) _T_2581;
  assign _T_2734 = _T_2692 & (* src = "crypto_accelerator.v:4835" *) _T_2557;
  assign _T_2736 = _T_2690 & (* src = "crypto_accelerator.v:4836" *) _T_2591;
  assign _T_2738 = _T_2700 & (* src = "crypto_accelerator.v:4837" *) _T_2562;
  assign _T_2740 = _T_2706 & (* src = "crypto_accelerator.v:4838" *) _T_2593;
  assign _T_2742 = _T_2698 & (* src = "crypto_accelerator.v:4839" *) _T_2560;
  assign _T_2897 = _T_2858 & (* src = "crypto_accelerator.v:4915" *) _T_2885;
  assign _T_2899 = _T_2833 & (* src = "crypto_accelerator.v:4916" *) _T_2849;
  assign _T_2903 = _T_2851 & (* src = "crypto_accelerator.v:4918" *) _T_2883;
  assign _T_2907 = _T_2860 & (* src = "crypto_accelerator.v:4920" *) _T_2887;
  assign _T_2909 = _T_2836 & (* src = "crypto_accelerator.v:4921" *) _T_2854;
  assign _T_2913 = _T_2870 & (* src = "crypto_accelerator.v:4923" *) _T_2868;
  assign _T_2917 = _T_2841 & (* src = "crypto_accelerator.v:4925" *) _T_2891;
  assign _T_2919 = _T_2872 & (* src = "crypto_accelerator.v:4926" *) _T_2889;
  assign _T_2923 = _T_2839 & (* src = "crypto_accelerator.v:4928" *) _T_2856;
  assign _T_2945 = _T_2939 & (* src = "crypto_accelerator.v:4939" *) _T_2935;
  assign _T_2953 = _T_2951 & (* src = "crypto_accelerator.v:4943" *) _T_2949;
  assign _T_2955 = _T_2947 & (* src = "crypto_accelerator.v:4944" *) _T_2943;
  assign _T_2957 = _T_2935 & (* src = "crypto_accelerator.v:4945" *) _T_2941;
  assign _T_2959 = _T_2949 & (* src = "crypto_accelerator.v:4946" *) _T_2957;
  assign _T_2963 = _T_2937 & (* src = "crypto_accelerator.v:4948" *) _T_2939;
  assign _T_2965 = _T_2943 & (* src = "crypto_accelerator.v:4949" *) _T_2963;
  assign _T_2987 = _T_2983 & (* src = "crypto_accelerator.v:4960" *) _T_2885;
  assign _T_2989 = _T_2975 & (* src = "crypto_accelerator.v:4961" *) _T_2849;
  assign _T_2991 = _T_2973 & (* src = "crypto_accelerator.v:4962" *) _T_2883;
  assign _T_2993 = _T_2981 & (* src = "crypto_accelerator.v:4963" *) _T_2887;
  assign _T_2995 = _T_2971 & (* src = "crypto_accelerator.v:4964" *) _T_2854;
  assign _T_2997 = _T_2969 & (* src = "crypto_accelerator.v:4965" *) _T_2868;
  assign _T_2999 = _T_2979 & (* src = "crypto_accelerator.v:4966" *) _T_2891;
  assign _T_3001 = _T_2985 & (* src = "crypto_accelerator.v:4967" *) _T_2889;
  assign _T_3003 = _T_2977 & (* src = "crypto_accelerator.v:4968" *) _T_2856;
  assign _T_3005 = _T_2983 & (* src = "crypto_accelerator.v:4969" *) _T_2858;
  assign _T_3007 = _T_2975 & (* src = "crypto_accelerator.v:4970" *) _T_2833;
  assign _T_3009 = _T_2973 & (* src = "crypto_accelerator.v:4971" *) _T_2851;
  assign _T_3011 = _T_2981 & (* src = "crypto_accelerator.v:4972" *) _T_2860;
  assign _T_3013 = _T_2971 & (* src = "crypto_accelerator.v:4973" *) _T_2836;
  assign _T_3015 = _T_2969 & (* src = "crypto_accelerator.v:4974" *) _T_2870;
  assign _T_3017 = _T_2979 & (* src = "crypto_accelerator.v:4975" *) _T_2841;
  assign _T_3019 = _T_2985 & (* src = "crypto_accelerator.v:4976" *) _T_2872;
  assign _T_3021 = _T_2977 & (* src = "crypto_accelerator.v:4977" *) _T_2839;
  assign _T_3176 = _T_3137 & (* src = "crypto_accelerator.v:5053" *) _T_3164;
  assign _T_3178 = _T_3112 & (* src = "crypto_accelerator.v:5054" *) _T_3128;
  assign _T_3182 = _T_3130 & (* src = "crypto_accelerator.v:5056" *) _T_3162;
  assign _T_3186 = _T_3139 & (* src = "crypto_accelerator.v:5058" *) _T_3166;
  assign _T_3188 = _T_3115 & (* src = "crypto_accelerator.v:5059" *) _T_3133;
  assign _T_3192 = _T_3149 & (* src = "crypto_accelerator.v:5061" *) _T_3147;
  assign _T_3196 = _T_3120 & (* src = "crypto_accelerator.v:5063" *) _T_3170;
  assign _T_3198 = _T_3151 & (* src = "crypto_accelerator.v:5064" *) _T_3168;
  assign _T_3202 = _T_3118 & (* src = "crypto_accelerator.v:5066" *) _T_3135;
  assign _T_3224 = _T_3218 & (* src = "crypto_accelerator.v:5077" *) _T_3214;
  assign _T_3232 = _T_3230 & (* src = "crypto_accelerator.v:5081" *) _T_3228;
  assign _T_3234 = _T_3226 & (* src = "crypto_accelerator.v:5082" *) _T_3222;
  assign _T_3236 = _T_3214 & (* src = "crypto_accelerator.v:5083" *) _T_3220;
  assign _T_3238 = _T_3228 & (* src = "crypto_accelerator.v:5084" *) _T_3236;
  assign _T_3242 = _T_3216 & (* src = "crypto_accelerator.v:5086" *) _T_3218;
  assign _T_3244 = _T_3222 & (* src = "crypto_accelerator.v:5087" *) _T_3242;
  assign _T_3266 = _T_3262 & (* src = "crypto_accelerator.v:5098" *) _T_3164;
  assign _T_3268 = _T_3254 & (* src = "crypto_accelerator.v:5099" *) _T_3128;
  assign _T_3270 = _T_3252 & (* src = "crypto_accelerator.v:5100" *) _T_3162;
  assign _T_3272 = _T_3260 & (* src = "crypto_accelerator.v:5101" *) _T_3166;
  assign _T_3274 = _T_3250 & (* src = "crypto_accelerator.v:5102" *) _T_3133;
  assign _T_3276 = _T_3248 & (* src = "crypto_accelerator.v:5103" *) _T_3147;
  assign _T_3278 = _T_3258 & (* src = "crypto_accelerator.v:5104" *) _T_3170;
  assign _T_3280 = _T_3264 & (* src = "crypto_accelerator.v:5105" *) _T_3168;
  assign _T_3282 = _T_3256 & (* src = "crypto_accelerator.v:5106" *) _T_3135;
  assign _T_3284 = _T_3262 & (* src = "crypto_accelerator.v:5107" *) _T_3137;
  assign _T_3286 = _T_3254 & (* src = "crypto_accelerator.v:5108" *) _T_3112;
  assign _T_3288 = _T_3252 & (* src = "crypto_accelerator.v:5109" *) _T_3130;
  assign _T_3290 = _T_3260 & (* src = "crypto_accelerator.v:5110" *) _T_3139;
  assign _T_3292 = _T_3250 & (* src = "crypto_accelerator.v:5111" *) _T_3115;
  assign _T_3294 = _T_3248 & (* src = "crypto_accelerator.v:5112" *) _T_3149;
  assign _T_3296 = _T_3258 & (* src = "crypto_accelerator.v:5113" *) _T_3120;
  assign _T_3298 = _T_3264 & (* src = "crypto_accelerator.v:5114" *) _T_3151;
  assign _T_3300 = _T_3256 & (* src = "crypto_accelerator.v:5115" *) _T_3118;
  assign _T_3456 = _T_3417 & (* src = "crypto_accelerator.v:5191" *) _T_3444;
  assign _T_3458 = _T_3392 & (* src = "crypto_accelerator.v:5192" *) _T_3408;
  assign _T_3462 = _T_3410 & (* src = "crypto_accelerator.v:5194" *) _T_3442;
  assign _T_3466 = _T_3419 & (* src = "crypto_accelerator.v:5196" *) _T_3446;
  assign _T_3468 = _T_3395 & (* src = "crypto_accelerator.v:5197" *) _T_3413;
  assign _T_3472 = _T_3429 & (* src = "crypto_accelerator.v:5199" *) _T_3427;
  assign _T_3476 = _T_3400 & (* src = "crypto_accelerator.v:5201" *) _T_3450;
  assign _T_3478 = _T_3431 & (* src = "crypto_accelerator.v:5202" *) _T_3448;
  assign _T_3482 = _T_3398 & (* src = "crypto_accelerator.v:5204" *) _T_3415;
  assign _T_3504 = _T_3498 & (* src = "crypto_accelerator.v:5215" *) _T_3494;
  assign _T_3512 = _T_3510 & (* src = "crypto_accelerator.v:5219" *) _T_3508;
  assign _T_3514 = _T_3506 & (* src = "crypto_accelerator.v:5220" *) _T_3502;
  assign _T_3516 = _T_3494 & (* src = "crypto_accelerator.v:5221" *) _T_3500;
  assign _T_3518 = _T_3508 & (* src = "crypto_accelerator.v:5222" *) _T_3516;
  assign _T_3522 = _T_3496 & (* src = "crypto_accelerator.v:5224" *) _T_3498;
  assign _T_3524 = _T_3502 & (* src = "crypto_accelerator.v:5225" *) _T_3522;
  assign _T_3546 = _T_3542 & (* src = "crypto_accelerator.v:5236" *) _T_3444;
  assign _T_3548 = _T_3534 & (* src = "crypto_accelerator.v:5237" *) _T_3408;
  assign _T_3550 = _T_3532 & (* src = "crypto_accelerator.v:5238" *) _T_3442;
  assign _T_3552 = _T_3540 & (* src = "crypto_accelerator.v:5239" *) _T_3446;
  assign _T_3554 = _T_3530 & (* src = "crypto_accelerator.v:5240" *) _T_3413;
  assign _T_3556 = _T_3528 & (* src = "crypto_accelerator.v:5241" *) _T_3427;
  assign _T_3558 = _T_3538 & (* src = "crypto_accelerator.v:5242" *) _T_3450;
  assign _T_3560 = _T_3544 & (* src = "crypto_accelerator.v:5243" *) _T_3448;
  assign _T_3562 = _T_3536 & (* src = "crypto_accelerator.v:5244" *) _T_3415;
  assign _T_3564 = _T_3542 & (* src = "crypto_accelerator.v:5245" *) _T_3417;
  assign _T_3566 = _T_3534 & (* src = "crypto_accelerator.v:5246" *) _T_3392;
  assign _T_3568 = _T_3532 & (* src = "crypto_accelerator.v:5247" *) _T_3410;
  assign _T_3570 = _T_3540 & (* src = "crypto_accelerator.v:5248" *) _T_3419;
  assign _T_3572 = _T_3530 & (* src = "crypto_accelerator.v:5249" *) _T_3395;
  assign _T_3574 = _T_3528 & (* src = "crypto_accelerator.v:5250" *) _T_3429;
  assign _T_3576 = _T_3538 & (* src = "crypto_accelerator.v:5251" *) _T_3400;
  assign _T_3578 = _T_3544 & (* src = "crypto_accelerator.v:5252" *) _T_3431;
  assign _T_3580 = _T_3536 & (* src = "crypto_accelerator.v:5253" *) _T_3398;
  assign _T_3735 = _T_3696 & (* src = "crypto_accelerator.v:5329" *) _T_3723;
  assign _T_3737 = _T_3671 & (* src = "crypto_accelerator.v:5330" *) _T_3687;
  assign _T_3741 = _T_3689 & (* src = "crypto_accelerator.v:5332" *) _T_3721;
  assign _T_3745 = _T_3698 & (* src = "crypto_accelerator.v:5334" *) _T_3725;
  assign _T_3747 = _T_3674 & (* src = "crypto_accelerator.v:5335" *) _T_3692;
  assign _T_3751 = _T_3708 & (* src = "crypto_accelerator.v:5337" *) _T_3706;
  assign _T_3755 = _T_3679 & (* src = "crypto_accelerator.v:5339" *) _T_3729;
  assign _T_3757 = _T_3710 & (* src = "crypto_accelerator.v:5340" *) _T_3727;
  assign _T_3761 = _T_3677 & (* src = "crypto_accelerator.v:5342" *) _T_3694;
  assign _T_3783 = _T_3777 & (* src = "crypto_accelerator.v:5353" *) _T_3773;
  assign _T_3791 = _T_3789 & (* src = "crypto_accelerator.v:5357" *) _T_3787;
  assign _T_3793 = _T_3785 & (* src = "crypto_accelerator.v:5358" *) _T_3781;
  assign _T_3795 = _T_3773 & (* src = "crypto_accelerator.v:5359" *) _T_3779;
  assign _T_3797 = _T_3787 & (* src = "crypto_accelerator.v:5360" *) _T_3795;
  assign _T_3801 = _T_3775 & (* src = "crypto_accelerator.v:5362" *) _T_3777;
  assign _T_3803 = _T_3781 & (* src = "crypto_accelerator.v:5363" *) _T_3801;
  assign _T_3825 = _T_3821 & (* src = "crypto_accelerator.v:5374" *) _T_3723;
  assign _T_3827 = _T_3813 & (* src = "crypto_accelerator.v:5375" *) _T_3687;
  assign _T_3829 = _T_3811 & (* src = "crypto_accelerator.v:5376" *) _T_3721;
  assign _T_3831 = _T_3819 & (* src = "crypto_accelerator.v:5377" *) _T_3725;
  assign _T_3833 = _T_3809 & (* src = "crypto_accelerator.v:5378" *) _T_3692;
  assign _T_3835 = _T_3807 & (* src = "crypto_accelerator.v:5379" *) _T_3706;
  assign _T_3837 = _T_3817 & (* src = "crypto_accelerator.v:5380" *) _T_3729;
  assign _T_3839 = _T_3823 & (* src = "crypto_accelerator.v:5381" *) _T_3727;
  assign _T_3841 = _T_3815 & (* src = "crypto_accelerator.v:5382" *) _T_3694;
  assign _T_3843 = _T_3821 & (* src = "crypto_accelerator.v:5383" *) _T_3696;
  assign _T_3845 = _T_3813 & (* src = "crypto_accelerator.v:5384" *) _T_3671;
  assign _T_3847 = _T_3811 & (* src = "crypto_accelerator.v:5385" *) _T_3689;
  assign _T_3849 = _T_3819 & (* src = "crypto_accelerator.v:5386" *) _T_3698;
  assign _T_3851 = _T_3809 & (* src = "crypto_accelerator.v:5387" *) _T_3674;
  assign _T_3853 = _T_3807 & (* src = "crypto_accelerator.v:5388" *) _T_3708;
  assign _T_3855 = _T_3817 & (* src = "crypto_accelerator.v:5389" *) _T_3679;
  assign _T_3857 = _T_3823 & (* src = "crypto_accelerator.v:5390" *) _T_3710;
  assign _T_3859 = _T_3815 & (* src = "crypto_accelerator.v:5391" *) _T_3677;
  assign _T_4014 = _T_3975 & (* src = "crypto_accelerator.v:5467" *) _T_4002;
  assign _T_4016 = _T_3950 & (* src = "crypto_accelerator.v:5468" *) _T_3966;
  assign _T_4020 = _T_3968 & (* src = "crypto_accelerator.v:5470" *) _T_4000;
  assign _T_4024 = _T_3977 & (* src = "crypto_accelerator.v:5472" *) _T_4004;
  assign _T_4026 = _T_3953 & (* src = "crypto_accelerator.v:5473" *) _T_3971;
  assign _T_4030 = _T_3987 & (* src = "crypto_accelerator.v:5475" *) _T_3985;
  assign _T_4034 = _T_3958 & (* src = "crypto_accelerator.v:5477" *) _T_4008;
  assign _T_4036 = _T_3989 & (* src = "crypto_accelerator.v:5478" *) _T_4006;
  assign _T_4040 = _T_3956 & (* src = "crypto_accelerator.v:5480" *) _T_3973;
  assign _T_4062 = _T_4056 & (* src = "crypto_accelerator.v:5491" *) _T_4052;
  assign _T_4070 = _T_4068 & (* src = "crypto_accelerator.v:5495" *) _T_4066;
  assign _T_4072 = _T_4064 & (* src = "crypto_accelerator.v:5496" *) _T_4060;
  assign _T_4074 = _T_4052 & (* src = "crypto_accelerator.v:5497" *) _T_4058;
  assign _T_4076 = _T_4066 & (* src = "crypto_accelerator.v:5498" *) _T_4074;
  assign _T_4080 = _T_4054 & (* src = "crypto_accelerator.v:5500" *) _T_4056;
  assign _T_4082 = _T_4060 & (* src = "crypto_accelerator.v:5501" *) _T_4080;
  assign _T_4104 = _T_4100 & (* src = "crypto_accelerator.v:5512" *) _T_4002;
  assign _T_4106 = _T_4092 & (* src = "crypto_accelerator.v:5513" *) _T_3966;
  assign _T_4108 = _T_4090 & (* src = "crypto_accelerator.v:5514" *) _T_4000;
  assign _T_4110 = _T_4098 & (* src = "crypto_accelerator.v:5515" *) _T_4004;
  assign _T_4112 = _T_4088 & (* src = "crypto_accelerator.v:5516" *) _T_3971;
  assign _T_4114 = _T_4086 & (* src = "crypto_accelerator.v:5517" *) _T_3985;
  assign _T_4116 = _T_4096 & (* src = "crypto_accelerator.v:5518" *) _T_4008;
  assign _T_4118 = _T_4102 & (* src = "crypto_accelerator.v:5519" *) _T_4006;
  assign _T_4120 = _T_4094 & (* src = "crypto_accelerator.v:5520" *) _T_3973;
  assign _T_4122 = _T_4100 & (* src = "crypto_accelerator.v:5521" *) _T_3975;
  assign _T_4124 = _T_4092 & (* src = "crypto_accelerator.v:5522" *) _T_3950;
  assign _T_4126 = _T_4090 & (* src = "crypto_accelerator.v:5523" *) _T_3968;
  assign _T_4128 = _T_4098 & (* src = "crypto_accelerator.v:5524" *) _T_3977;
  assign _T_4130 = _T_4088 & (* src = "crypto_accelerator.v:5525" *) _T_3953;
  assign _T_4132 = _T_4086 & (* src = "crypto_accelerator.v:5526" *) _T_3987;
  assign _T_4134 = _T_4096 & (* src = "crypto_accelerator.v:5527" *) _T_3958;
  assign _T_4136 = _T_4102 & (* src = "crypto_accelerator.v:5528" *) _T_3989;
  assign _T_4138 = _T_4094 & (* src = "crypto_accelerator.v:5529" *) _T_3956;
  assign _T_4293 = _T_4254 & (* src = "crypto_accelerator.v:5605" *) _T_4281;
  assign _T_4295 = _T_4229 & (* src = "crypto_accelerator.v:5606" *) _T_4245;
  assign _T_4299 = _T_4247 & (* src = "crypto_accelerator.v:5608" *) _T_4279;
  assign _T_4303 = _T_4256 & (* src = "crypto_accelerator.v:5610" *) _T_4283;
  assign _T_4305 = _T_4232 & (* src = "crypto_accelerator.v:5611" *) _T_4250;
  assign _T_4309 = _T_4266 & (* src = "crypto_accelerator.v:5613" *) _T_4264;
  assign _T_4313 = _T_4237 & (* src = "crypto_accelerator.v:5615" *) _T_4287;
  assign _T_4315 = _T_4268 & (* src = "crypto_accelerator.v:5616" *) _T_4285;
  assign _T_4319 = _T_4235 & (* src = "crypto_accelerator.v:5618" *) _T_4252;
  assign _T_4341 = _T_4335 & (* src = "crypto_accelerator.v:5629" *) _T_4331;
  assign _T_4349 = _T_4347 & (* src = "crypto_accelerator.v:5633" *) _T_4345;
  assign _T_4351 = _T_4343 & (* src = "crypto_accelerator.v:5634" *) _T_4339;
  assign _T_4353 = _T_4331 & (* src = "crypto_accelerator.v:5635" *) _T_4337;
  assign _T_4355 = _T_4345 & (* src = "crypto_accelerator.v:5636" *) _T_4353;
  assign _T_4359 = _T_4333 & (* src = "crypto_accelerator.v:5638" *) _T_4335;
  assign _T_4361 = _T_4339 & (* src = "crypto_accelerator.v:5639" *) _T_4359;
  assign _T_4383 = _T_4379 & (* src = "crypto_accelerator.v:5650" *) _T_4281;
  assign _T_4385 = _T_4371 & (* src = "crypto_accelerator.v:5651" *) _T_4245;
  assign _T_4387 = _T_4369 & (* src = "crypto_accelerator.v:5652" *) _T_4279;
  assign _T_4389 = _T_4377 & (* src = "crypto_accelerator.v:5653" *) _T_4283;
  assign _T_4391 = _T_4367 & (* src = "crypto_accelerator.v:5654" *) _T_4250;
  assign _T_4393 = _T_4365 & (* src = "crypto_accelerator.v:5655" *) _T_4264;
  assign _T_4395 = _T_4375 & (* src = "crypto_accelerator.v:5656" *) _T_4287;
  assign _T_4397 = _T_4381 & (* src = "crypto_accelerator.v:5657" *) _T_4285;
  assign _T_4399 = _T_4373 & (* src = "crypto_accelerator.v:5658" *) _T_4252;
  assign _T_4401 = _T_4379 & (* src = "crypto_accelerator.v:5659" *) _T_4254;
  assign _T_4403 = _T_4371 & (* src = "crypto_accelerator.v:5660" *) _T_4229;
  assign _T_4405 = _T_4369 & (* src = "crypto_accelerator.v:5661" *) _T_4247;
  assign _T_4407 = _T_4377 & (* src = "crypto_accelerator.v:5662" *) _T_4256;
  assign _T_4409 = _T_4367 & (* src = "crypto_accelerator.v:5663" *) _T_4232;
  assign _T_4411 = _T_4365 & (* src = "crypto_accelerator.v:5664" *) _T_4266;
  assign _T_4413 = _T_4375 & (* src = "crypto_accelerator.v:5665" *) _T_4237;
  assign _T_4415 = _T_4381 & (* src = "crypto_accelerator.v:5666" *) _T_4268;
  assign _T_4417 = _T_4373 & (* src = "crypto_accelerator.v:5667" *) _T_4235;
  assign _T_4535 = _T_4534 & (* src = "crypto_accelerator.v:5948" *) 8'b10000000;
  assign _T_4539 = _T_4538 & (* src = "crypto_accelerator.v:5952" *) 8'b11111111;
  assign _T_4542 = _T_4541 & (* src = "crypto_accelerator.v:5954" *) 8'b10000000;
  assign _T_4546 = _T_4545 & (* src = "crypto_accelerator.v:5958" *) 8'b11111111;
  assign _T_4550 = _T_4549 & (* src = "crypto_accelerator.v:5961" *) 8'b10000000;
  assign _T_4554 = _T_4553 & (* src = "crypto_accelerator.v:5965" *) 8'b11111111;
  assign _T_4557 = _T_4556 & (* src = "crypto_accelerator.v:5967" *) 8'b10000000;
  assign _T_4561 = _T_4560 & (* src = "crypto_accelerator.v:5971" *) 8'b11111111;
  assign _T_4569 = _T_4568 & (* src = "crypto_accelerator.v:5982" *) 8'b10000000;
  assign _T_4573 = _T_4572 & (* src = "crypto_accelerator.v:5986" *) 8'b11111111;
  assign _T_4576 = _T_4575 & (* src = "crypto_accelerator.v:5988" *) 8'b10000000;
  assign _T_4580 = _T_4579 & (* src = "crypto_accelerator.v:5992" *) 8'b11111111;
  assign _T_4584 = _T_4583 & (* src = "crypto_accelerator.v:5995" *) 8'b10000000;
  assign _T_4588 = _T_4587 & (* src = "crypto_accelerator.v:5999" *) 8'b11111111;
  assign _T_4591 = _T_4590 & (* src = "crypto_accelerator.v:6001" *) 8'b10000000;
  assign _T_4595[7:0] = _T_4594 & (* src = "crypto_accelerator.v:6005" *) 8'b11111111;
  assign _T_4603 = _T_4602 & (* src = "crypto_accelerator.v:6016" *) 8'b10000000;
  assign _T_4607 = _T_4606 & (* src = "crypto_accelerator.v:6020" *) 8'b11111111;
  assign _T_4610 = _T_4609 & (* src = "crypto_accelerator.v:6022" *) 8'b10000000;
  assign _T_4614 = _T_4613 & (* src = "crypto_accelerator.v:6026" *) 8'b11111111;
  assign _T_4618 = _T_4617 & (* src = "crypto_accelerator.v:6029" *) 8'b10000000;
  assign _T_4622 = _T_4621 & (* src = "crypto_accelerator.v:6033" *) 8'b11111111;
  assign _T_4625 = _T_4624 & (* src = "crypto_accelerator.v:6035" *) 8'b10000000;
  assign _T_4629[7:0] = _T_4628 & (* src = "crypto_accelerator.v:6039" *) 8'b11111111;
  assign _T_4637 = _T_4636 & (* src = "crypto_accelerator.v:6050" *) 8'b10000000;
  assign _T_4641 = _T_4640 & (* src = "crypto_accelerator.v:6054" *) 8'b11111111;
  assign _T_4644 = _T_4643 & (* src = "crypto_accelerator.v:6056" *) 8'b10000000;
  assign _T_4648 = _T_4647 & (* src = "crypto_accelerator.v:6060" *) 8'b11111111;
  assign _T_4652 = _T_4651 & (* src = "crypto_accelerator.v:6063" *) 8'b10000000;
  assign _T_4656 = _T_4655 & (* src = "crypto_accelerator.v:6067" *) 8'b11111111;
  assign _T_4659 = _T_4658 & (* src = "crypto_accelerator.v:6069" *) 8'b10000000;
  assign _T_4663[7:0] = _T_4662 & (* src = "crypto_accelerator.v:6073" *) 8'b11111111;
  assign _T_4747 = io_ready & (* src = "crypto_accelerator.v:6102" *) io_dataValid;
  assign io_shift = _T_4770 & (* src = "crypto_accelerator.v:6148" *) _GEN_292;
  assign _T = ! (* src = "crypto_accelerator.v:3477" *) state;
  assign _T_1 = state == (* src = "crypto_accelerator.v:3478" *) 5'b11110;
  assign _0018_ = ! (* src = "crypto_accelerator.v:5819" *) keyEndAddr;
  assign _0019_ = 3'b001 == (* src = "crypto_accelerator.v:5835" *) keyEndAddr;
  assign _0020_ = 3'b010 == (* src = "crypto_accelerator.v:5851" *) keyEndAddr;
  assign _0021_ = 3'b011 == (* src = "crypto_accelerator.v:5867" *) keyEndAddr;
  assign _0022_ = 3'b100 == (* src = "crypto_accelerator.v:5883" *) keyEndAddr;
  assign _0023_ = 3'b101 == (* src = "crypto_accelerator.v:5899" *) keyEndAddr;
  assign _0024_ = 3'b110 == (* src = "crypto_accelerator.v:5915" *) keyEndAddr;
  assign _T_4771 = state == (* src = "crypto_accelerator.v:6105" *) 1'b1;
  assign _T_4775 = state == (* src = "crypto_accelerator.v:6108" *) { 1'b1, _GEN_327 };
  assign _T_4536 = | (* src = "crypto_accelerator.v:5949" *) _T_4535;
  assign _T_4543 = | (* src = "crypto_accelerator.v:5955" *) _T_4542;
  assign _T_4551 = | (* src = "crypto_accelerator.v:5962" *) _T_4550;
  assign _T_4558 = | (* src = "crypto_accelerator.v:5968" *) _T_4557;
  assign _T_4570 = | (* src = "crypto_accelerator.v:5983" *) _T_4569;
  assign _T_4577 = | (* src = "crypto_accelerator.v:5989" *) _T_4576;
  assign _T_4585 = | (* src = "crypto_accelerator.v:5996" *) _T_4584;
  assign _T_4592 = | (* src = "crypto_accelerator.v:6002" *) _T_4591;
  assign _T_4604 = | (* src = "crypto_accelerator.v:6017" *) _T_4603;
  assign _T_4611 = | (* src = "crypto_accelerator.v:6023" *) _T_4610;
  assign _T_4619 = | (* src = "crypto_accelerator.v:6030" *) _T_4618;
  assign _T_4626 = | (* src = "crypto_accelerator.v:6036" *) _T_4625;
  assign _T_4638 = | (* src = "crypto_accelerator.v:6051" *) _T_4637;
  assign _T_4645 = | (* src = "crypto_accelerator.v:6057" *) _T_4644;
  assign _T_4653 = | (* src = "crypto_accelerator.v:6064" *) _T_4652;
  assign _T_4660 = | (* src = "crypto_accelerator.v:6070" *) _T_4659;
  assign _T_44 = ~ (* src = "crypto_accelerator.v:3500" *) _T_43;
  assign _T_47 = ~ (* src = "crypto_accelerator.v:3502" *) _T_46;
  assign _T_52 = ~ (* src = "crypto_accelerator.v:3505" *) _T_51;
  assign _T_57 = ~ (* src = "crypto_accelerator.v:3508" *) _T_56;
  assign _T_62 = ~ (* src = "crypto_accelerator.v:3511" *) _T_61;
  assign _T_71 = ~ (* src = "crypto_accelerator.v:3516" *) _T_70;
  assign _T_76 = ~ (* src = "crypto_accelerator.v:3519" *) _T_75;
  assign _T_83 = ~ (* src = "crypto_accelerator.v:3523" *) _T_82;
  assign _T_86 = ~ (* src = "crypto_accelerator.v:3525" *) _T_85;
  assign _T_89 = ~ (* src = "crypto_accelerator.v:3527" *) _T_88;
  assign _T_323 = ~ (* src = "crypto_accelerator.v:3638" *) _T_322;
  assign _T_326 = ~ (* src = "crypto_accelerator.v:3640" *) _T_325;
  assign _T_331 = ~ (* src = "crypto_accelerator.v:3643" *) _T_330;
  assign _T_336 = ~ (* src = "crypto_accelerator.v:3646" *) _T_335;
  assign _T_341 = ~ (* src = "crypto_accelerator.v:3649" *) _T_340;
  assign _T_350 = ~ (* src = "crypto_accelerator.v:3654" *) _T_349;
  assign _T_355 = ~ (* src = "crypto_accelerator.v:3657" *) _T_354;
  assign _T_362 = ~ (* src = "crypto_accelerator.v:3661" *) _T_361;
  assign _T_365 = ~ (* src = "crypto_accelerator.v:3663" *) _T_364;
  assign _T_368 = ~ (* src = "crypto_accelerator.v:3665" *) _T_367;
  assign _T_602 = ~ (* src = "crypto_accelerator.v:3776" *) _T_601;
  assign _T_605 = ~ (* src = "crypto_accelerator.v:3778" *) _T_604;
  assign _T_610 = ~ (* src = "crypto_accelerator.v:3781" *) _T_609;
  assign _T_615 = ~ (* src = "crypto_accelerator.v:3784" *) _T_614;
  assign _T_620 = ~ (* src = "crypto_accelerator.v:3787" *) _T_619;
  assign _T_629 = ~ (* src = "crypto_accelerator.v:3792" *) _T_628;
  assign _T_634 = ~ (* src = "crypto_accelerator.v:3795" *) _T_633;
  assign _T_641 = ~ (* src = "crypto_accelerator.v:3799" *) _T_640;
  assign _T_644 = ~ (* src = "crypto_accelerator.v:3801" *) _T_643;
  assign _T_647 = ~ (* src = "crypto_accelerator.v:3803" *) _T_646;
  assign _T_881 = ~ (* src = "crypto_accelerator.v:3914" *) _T_880;
  assign _T_884 = ~ (* src = "crypto_accelerator.v:3916" *) _T_883;
  assign _T_889 = ~ (* src = "crypto_accelerator.v:3919" *) _T_888;
  assign _T_894 = ~ (* src = "crypto_accelerator.v:3922" *) _T_893;
  assign _T_899 = ~ (* src = "crypto_accelerator.v:3925" *) _T_898;
  assign _T_908 = ~ (* src = "crypto_accelerator.v:3930" *) _T_907;
  assign _T_913 = ~ (* src = "crypto_accelerator.v:3933" *) _T_912;
  assign _T_920 = ~ (* src = "crypto_accelerator.v:3937" *) _T_919;
  assign _T_923 = ~ (* src = "crypto_accelerator.v:3939" *) _T_922;
  assign _T_926 = ~ (* src = "crypto_accelerator.v:3941" *) _T_925;
  assign _T_1161 = ~ (* src = "crypto_accelerator.v:4052" *) _T_1160;
  assign _T_1164 = ~ (* src = "crypto_accelerator.v:4054" *) _T_1163;
  assign _T_1169 = ~ (* src = "crypto_accelerator.v:4057" *) _T_1168;
  assign _T_1174 = ~ (* src = "crypto_accelerator.v:4060" *) _T_1173;
  assign _T_1179 = ~ (* src = "crypto_accelerator.v:4063" *) _T_1178;
  assign _T_1188 = ~ (* src = "crypto_accelerator.v:4068" *) _T_1187;
  assign _T_1193 = ~ (* src = "crypto_accelerator.v:4071" *) _T_1192;
  assign _T_1200 = ~ (* src = "crypto_accelerator.v:4075" *) _T_1199;
  assign _T_1203 = ~ (* src = "crypto_accelerator.v:4077" *) _T_1202;
  assign _T_1206 = ~ (* src = "crypto_accelerator.v:4079" *) _T_1205;
  assign _T_1440 = ~ (* src = "crypto_accelerator.v:4190" *) _T_1439;
  assign _T_1443 = ~ (* src = "crypto_accelerator.v:4192" *) _T_1442;
  assign _T_1448 = ~ (* src = "crypto_accelerator.v:4195" *) _T_1447;
  assign _T_1453 = ~ (* src = "crypto_accelerator.v:4198" *) _T_1452;
  assign _T_1458 = ~ (* src = "crypto_accelerator.v:4201" *) _T_1457;
  assign _T_1467 = ~ (* src = "crypto_accelerator.v:4206" *) _T_1466;
  assign _T_1472 = ~ (* src = "crypto_accelerator.v:4209" *) _T_1471;
  assign _T_1479 = ~ (* src = "crypto_accelerator.v:4213" *) _T_1478;
  assign _T_1482 = ~ (* src = "crypto_accelerator.v:4215" *) _T_1481;
  assign _T_1485 = ~ (* src = "crypto_accelerator.v:4217" *) _T_1484;
  assign _T_1719 = ~ (* src = "crypto_accelerator.v:4328" *) _T_1718;
  assign _T_1722 = ~ (* src = "crypto_accelerator.v:4330" *) _T_1721;
  assign _T_1727 = ~ (* src = "crypto_accelerator.v:4333" *) _T_1726;
  assign _T_1732 = ~ (* src = "crypto_accelerator.v:4336" *) _T_1731;
  assign _T_1737 = ~ (* src = "crypto_accelerator.v:4339" *) _T_1736;
  assign _T_1746 = ~ (* src = "crypto_accelerator.v:4344" *) _T_1745;
  assign _T_1751 = ~ (* src = "crypto_accelerator.v:4347" *) _T_1750;
  assign _T_1758 = ~ (* src = "crypto_accelerator.v:4351" *) _T_1757;
  assign _T_1761 = ~ (* src = "crypto_accelerator.v:4353" *) _T_1760;
  assign _T_1764 = ~ (* src = "crypto_accelerator.v:4355" *) _T_1763;
  assign _T_1998 = ~ (* src = "crypto_accelerator.v:4466" *) _T_1997;
  assign _T_2001 = ~ (* src = "crypto_accelerator.v:4468" *) _T_2000;
  assign _T_2006 = ~ (* src = "crypto_accelerator.v:4471" *) _T_2005;
  assign _T_2011 = ~ (* src = "crypto_accelerator.v:4474" *) _T_2010;
  assign _T_2016 = ~ (* src = "crypto_accelerator.v:4477" *) _T_2015;
  assign _T_2025 = ~ (* src = "crypto_accelerator.v:4482" *) _T_2024;
  assign _T_2030 = ~ (* src = "crypto_accelerator.v:4485" *) _T_2029;
  assign _T_2037 = ~ (* src = "crypto_accelerator.v:4489" *) _T_2036;
  assign _T_2040 = ~ (* src = "crypto_accelerator.v:4491" *) _T_2039;
  assign _T_2043 = ~ (* src = "crypto_accelerator.v:4493" *) _T_2042;
  assign _T_2278 = ~ (* src = "crypto_accelerator.v:4604" *) _T_2277;
  assign _T_2281 = ~ (* src = "crypto_accelerator.v:4606" *) _T_2280;
  assign _T_2286 = ~ (* src = "crypto_accelerator.v:4609" *) _T_2285;
  assign _T_2291 = ~ (* src = "crypto_accelerator.v:4612" *) _T_2290;
  assign _T_2296 = ~ (* src = "crypto_accelerator.v:4615" *) _T_2295;
  assign _T_2305 = ~ (* src = "crypto_accelerator.v:4620" *) _T_2304;
  assign _T_2310 = ~ (* src = "crypto_accelerator.v:4623" *) _T_2309;
  assign _T_2317 = ~ (* src = "crypto_accelerator.v:4627" *) _T_2316;
  assign _T_2320 = ~ (* src = "crypto_accelerator.v:4629" *) _T_2319;
  assign _T_2323 = ~ (* src = "crypto_accelerator.v:4631" *) _T_2322;
  assign _T_2557 = ~ (* src = "crypto_accelerator.v:4742" *) _T_2556;
  assign _T_2560 = ~ (* src = "crypto_accelerator.v:4744" *) _T_2559;
  assign _T_2565 = ~ (* src = "crypto_accelerator.v:4747" *) _T_2564;
  assign _T_2570 = ~ (* src = "crypto_accelerator.v:4750" *) _T_2569;
  assign _T_2575 = ~ (* src = "crypto_accelerator.v:4753" *) _T_2574;
  assign _T_2584 = ~ (* src = "crypto_accelerator.v:4758" *) _T_2583;
  assign _T_2589 = ~ (* src = "crypto_accelerator.v:4761" *) _T_2588;
  assign _T_2596 = ~ (* src = "crypto_accelerator.v:4765" *) _T_2595;
  assign _T_2599 = ~ (* src = "crypto_accelerator.v:4767" *) _T_2598;
  assign _T_2602 = ~ (* src = "crypto_accelerator.v:4769" *) _T_2601;
  assign _T_2836 = ~ (* src = "crypto_accelerator.v:4880" *) _T_2835;
  assign _T_2839 = ~ (* src = "crypto_accelerator.v:4882" *) _T_2838;
  assign _T_2844 = ~ (* src = "crypto_accelerator.v:4885" *) _T_2843;
  assign _T_2849 = ~ (* src = "crypto_accelerator.v:4888" *) _T_2848;
  assign _T_2854 = ~ (* src = "crypto_accelerator.v:4891" *) _T_2853;
  assign _T_2863 = ~ (* src = "crypto_accelerator.v:4896" *) _T_2862;
  assign _T_2868 = ~ (* src = "crypto_accelerator.v:4899" *) _T_2867;
  assign _T_2875 = ~ (* src = "crypto_accelerator.v:4903" *) _T_2874;
  assign _T_2878 = ~ (* src = "crypto_accelerator.v:4905" *) _T_2877;
  assign _T_2881 = ~ (* src = "crypto_accelerator.v:4907" *) _T_2880;
  assign _T_3115 = ~ (* src = "crypto_accelerator.v:5018" *) _T_3114;
  assign _T_3118 = ~ (* src = "crypto_accelerator.v:5020" *) _T_3117;
  assign _T_3123 = ~ (* src = "crypto_accelerator.v:5023" *) _T_3122;
  assign _T_3128 = ~ (* src = "crypto_accelerator.v:5026" *) _T_3127;
  assign _T_3133 = ~ (* src = "crypto_accelerator.v:5029" *) _T_3132;
  assign _T_3142 = ~ (* src = "crypto_accelerator.v:5034" *) _T_3141;
  assign _T_3147 = ~ (* src = "crypto_accelerator.v:5037" *) _T_3146;
  assign _T_3154 = ~ (* src = "crypto_accelerator.v:5041" *) _T_3153;
  assign _T_3157 = ~ (* src = "crypto_accelerator.v:5043" *) _T_3156;
  assign _T_3160 = ~ (* src = "crypto_accelerator.v:5045" *) _T_3159;
  assign _T_3395 = ~ (* src = "crypto_accelerator.v:5156" *) _T_3394;
  assign _T_3398 = ~ (* src = "crypto_accelerator.v:5158" *) _T_3397;
  assign _T_3403 = ~ (* src = "crypto_accelerator.v:5161" *) _T_3402;
  assign _T_3408 = ~ (* src = "crypto_accelerator.v:5164" *) _T_3407;
  assign _T_3413 = ~ (* src = "crypto_accelerator.v:5167" *) _T_3412;
  assign _T_3422 = ~ (* src = "crypto_accelerator.v:5172" *) _T_3421;
  assign _T_3427 = ~ (* src = "crypto_accelerator.v:5175" *) _T_3426;
  assign _T_3434 = ~ (* src = "crypto_accelerator.v:5179" *) _T_3433;
  assign _T_3437 = ~ (* src = "crypto_accelerator.v:5181" *) _T_3436;
  assign _T_3440 = ~ (* src = "crypto_accelerator.v:5183" *) _T_3439;
  assign _T_3674 = ~ (* src = "crypto_accelerator.v:5294" *) _T_3673;
  assign _T_3677 = ~ (* src = "crypto_accelerator.v:5296" *) _T_3676;
  assign _T_3682 = ~ (* src = "crypto_accelerator.v:5299" *) _T_3681;
  assign _T_3687 = ~ (* src = "crypto_accelerator.v:5302" *) _T_3686;
  assign _T_3692 = ~ (* src = "crypto_accelerator.v:5305" *) _T_3691;
  assign _T_3701 = ~ (* src = "crypto_accelerator.v:5310" *) _T_3700;
  assign _T_3706 = ~ (* src = "crypto_accelerator.v:5313" *) _T_3705;
  assign _T_3713 = ~ (* src = "crypto_accelerator.v:5317" *) _T_3712;
  assign _T_3716 = ~ (* src = "crypto_accelerator.v:5319" *) _T_3715;
  assign _T_3719 = ~ (* src = "crypto_accelerator.v:5321" *) _T_3718;
  assign _T_3953 = ~ (* src = "crypto_accelerator.v:5432" *) _T_3952;
  assign _T_3956 = ~ (* src = "crypto_accelerator.v:5434" *) _T_3955;
  assign _T_3961 = ~ (* src = "crypto_accelerator.v:5437" *) _T_3960;
  assign _T_3966 = ~ (* src = "crypto_accelerator.v:5440" *) _T_3965;
  assign _T_3971 = ~ (* src = "crypto_accelerator.v:5443" *) _T_3970;
  assign _T_3980 = ~ (* src = "crypto_accelerator.v:5448" *) _T_3979;
  assign _T_3985 = ~ (* src = "crypto_accelerator.v:5451" *) _T_3984;
  assign _T_3992 = ~ (* src = "crypto_accelerator.v:5455" *) _T_3991;
  assign _T_3995 = ~ (* src = "crypto_accelerator.v:5457" *) _T_3994;
  assign _T_3998 = ~ (* src = "crypto_accelerator.v:5459" *) _T_3997;
  assign _T_4232 = ~ (* src = "crypto_accelerator.v:5570" *) _T_4231;
  assign _T_4235 = ~ (* src = "crypto_accelerator.v:5572" *) _T_4234;
  assign _T_4240 = ~ (* src = "crypto_accelerator.v:5575" *) _T_4239;
  assign _T_4245 = ~ (* src = "crypto_accelerator.v:5578" *) _T_4244;
  assign _T_4250 = ~ (* src = "crypto_accelerator.v:5581" *) _T_4249;
  assign _T_4259 = ~ (* src = "crypto_accelerator.v:5586" *) _T_4258;
  assign _T_4264 = ~ (* src = "crypto_accelerator.v:5589" *) _T_4263;
  assign _T_4271 = ~ (* src = "crypto_accelerator.v:5593" *) _T_4270;
  assign _T_4274 = ~ (* src = "crypto_accelerator.v:5595" *) _T_4273;
  assign _T_4277 = ~ (* src = "crypto_accelerator.v:5597" *) _T_4276;
  assign _T_4770 = ~ (* src = "crypto_accelerator.v:6104" *) io_ready;
  assign _GEN_292 = _T_4771 | (* src = "crypto_accelerator.v:6110" *) state[0];
  assign io_ready = _T | (* src = "crypto_accelerator.v:6149" *) _T_1;
  always @(posedge clock)
      state <= _0017_;
  always @(posedge clock)
      matrix_0_0 <= _0001_;
  always @(posedge clock)
      matrix_0_1 <= _0002_;
  always @(posedge clock)
      matrix_0_2 <= _0003_;
  always @(posedge clock)
      matrix_0_3 <= _0004_;
  always @(posedge clock)
      matrix_1_0 <= _0005_;
  always @(posedge clock)
      matrix_1_1 <= _0006_;
  always @(posedge clock)
      matrix_1_2 <= _0007_;
  always @(posedge clock)
      matrix_1_3 <= _0008_;
  always @(posedge clock)
      matrix_2_0 <= _0009_;
  always @(posedge clock)
      matrix_2_1 <= _0010_;
  always @(posedge clock)
      matrix_2_2 <= _0011_;
  always @(posedge clock)
      matrix_2_3 <= _0012_;
  always @(posedge clock)
      matrix_3_0 <= _0013_;
  always @(posedge clock)
      matrix_3_1 <= _0014_;
  always @(posedge clock)
      matrix_3_2 <= _0015_;
  always @(posedge clock)
      matrix_3_3 <= _0016_;
  always @(posedge clock)
      ctSaved <= _0000_;
  assign _0000_ = _T_4747 ? (* src = "crypto_accelerator.v:6255" *) io_dataIn : ctSaved;
  assign _0025_ = _T_4747 ? (* src = "crypto_accelerator.v:6463" *) io_dataIn[7:0] : matrix_3_3;
  assign _0026_ = _T_4775 ? (* src = "crypto_accelerator.v:6458" *) xorOut_3_3 : MixColsModule_io_out_3_3;
  assign _0027_ = state[0] ? (* src = "crypto_accelerator.v:6456" *) _0026_ : { _T_4476, _T_4477, _T_4478, _T_4479, _T_4480, _T_4481, _T_4482, _T_4483 };
  assign _0028_ = _T_4771 ? (* src = "crypto_accelerator.v:6454" *) _T_4726[7:0] : _0027_;
  assign _0016_ = io_ready ? (* src = "crypto_accelerator.v:6453" *) _0025_ : _0028_;
  assign _0029_ = _T_4747 ? (* src = "crypto_accelerator.v:6450" *) io_dataIn[15:8] : matrix_3_2;
  assign _0030_ = _T_4775 ? (* src = "crypto_accelerator.v:6445" *) xorOut_3_2 : MixColsModule_io_out_3_2;
  assign _0031_ = state[0] ? (* src = "crypto_accelerator.v:6443" *) _0030_ : { _T_4197, _T_4198, _T_4199, _T_4200, _T_4201, _T_4202, _T_4203, _T_4204 };
  assign _0032_ = _T_4771 ? (* src = "crypto_accelerator.v:6441" *) _T_4726[15:8] : _0031_;
  assign _0015_ = io_ready ? (* src = "crypto_accelerator.v:6440" *) _0029_ : _0032_;
  assign _0033_ = _T_4747 ? (* src = "crypto_accelerator.v:6437" *) io_dataIn[23:16] : matrix_3_1;
  assign _0034_ = _T_4775 ? (* src = "crypto_accelerator.v:6432" *) xorOut_3_1 : MixColsModule_io_out_3_1;
  assign _0035_ = state[0] ? (* src = "crypto_accelerator.v:6430" *) _0034_ : { _T_3918, _T_3919, _T_3920, _T_3921, _T_3922, _T_3923, _T_3924, _T_3925 };
  assign _0036_ = _T_4771 ? (* src = "crypto_accelerator.v:6428" *) _T_4726[23:16] : _0035_;
  assign _0014_ = io_ready ? (* src = "crypto_accelerator.v:6427" *) _0033_ : _0036_;
  assign _0037_ = _T_4747 ? (* src = "crypto_accelerator.v:6424" *) io_dataIn[31:24] : matrix_3_0;
  assign _0038_ = _T_4775 ? (* src = "crypto_accelerator.v:6419" *) xorOut_3_0 : MixColsModule_io_out_3_0;
  assign _0039_ = state[0] ? (* src = "crypto_accelerator.v:6417" *) _0038_ : { _T_3639, _T_3640, _T_3641, _T_3642, _T_3643, _T_3644, _T_3645, _T_3646 };
  assign _0040_ = _T_4771 ? (* src = "crypto_accelerator.v:6415" *) _T_4726[31:24] : _0039_;
  assign _0013_ = io_ready ? (* src = "crypto_accelerator.v:6414" *) _0037_ : _0040_;
  assign _0041_ = _T_4747 ? (* src = "crypto_accelerator.v:6411" *) io_dataIn[39:32] : matrix_2_3;
  assign _0042_ = _T_4775 ? (* src = "crypto_accelerator.v:6406" *) xorOut_2_3 : MixColsModule_io_out_2_3;
  assign _0043_ = state[0] ? (* src = "crypto_accelerator.v:6404" *) _0042_ : { _T_3359, _T_3360, _T_3361, _T_3362, _T_3363, _T_3364, _T_3365, _T_3366 };
  assign _0044_ = _T_4771 ? (* src = "crypto_accelerator.v:6402" *) _T_4726[39:32] : _0043_;
  assign _0012_ = io_ready ? (* src = "crypto_accelerator.v:6401" *) _0041_ : _0044_;
  assign _0045_ = _T_4747 ? (* src = "crypto_accelerator.v:6398" *) io_dataIn[47:40] : matrix_2_2;
  assign _0046_ = _T_4775 ? (* src = "crypto_accelerator.v:6393" *) xorOut_2_2 : MixColsModule_io_out_2_2;
  assign _0047_ = state[0] ? (* src = "crypto_accelerator.v:6391" *) _0046_ : { _T_3080, _T_3081, _T_3082, _T_3083, _T_3084, _T_3085, _T_3086, _T_3087 };
  assign _0048_ = _T_4771 ? (* src = "crypto_accelerator.v:6389" *) _T_4726[47:40] : _0047_;
  assign _0011_ = io_ready ? (* src = "crypto_accelerator.v:6388" *) _0045_ : _0048_;
  assign _0049_ = _T_4747 ? (* src = "crypto_accelerator.v:6385" *) io_dataIn[55:48] : matrix_2_1;
  assign _0050_ = _T_4775 ? (* src = "crypto_accelerator.v:6380" *) xorOut_2_1 : MixColsModule_io_out_2_1;
  assign _0051_ = state[0] ? (* src = "crypto_accelerator.v:6378" *) _0050_ : { _T_2801, _T_2802, _T_2803, _T_2804, _T_2805, _T_2806, _T_2807, _T_2808 };
  assign _0052_ = _T_4771 ? (* src = "crypto_accelerator.v:6376" *) _T_4726[55:48] : _0051_;
  assign _0010_ = io_ready ? (* src = "crypto_accelerator.v:6375" *) _0049_ : _0052_;
  assign _0053_ = _T_4747 ? (* src = "crypto_accelerator.v:6372" *) io_dataIn[63:56] : matrix_2_0;
  assign _0054_ = _T_4775 ? (* src = "crypto_accelerator.v:6367" *) xorOut_2_0 : MixColsModule_io_out_2_0;
  assign _0055_ = state[0] ? (* src = "crypto_accelerator.v:6365" *) _0054_ : { _T_2522, _T_2523, _T_2524, _T_2525, _T_2526, _T_2527, _T_2528, _T_2529 };
  assign _0056_ = _T_4771 ? (* src = "crypto_accelerator.v:6363" *) _T_4726[63:56] : _0055_;
  assign _0009_ = io_ready ? (* src = "crypto_accelerator.v:6362" *) _0053_ : _0056_;
  assign _0057_ = _T_4747 ? (* src = "crypto_accelerator.v:6359" *) io_dataIn[71:64] : matrix_1_3;
  assign _0058_ = _T_4775 ? (* src = "crypto_accelerator.v:6354" *) xorOut_1_3 : MixColsModule_io_out_1_3;
  assign _0059_ = state[0] ? (* src = "crypto_accelerator.v:6352" *) _0058_ : { _T_2242, _T_2243, _T_2244, _T_2245, _T_2246, _T_2247, _T_2248, _T_2249 };
  assign _0060_ = _T_4771 ? (* src = "crypto_accelerator.v:6350" *) _T_4726[71:64] : _0059_;
  assign _0008_ = io_ready ? (* src = "crypto_accelerator.v:6349" *) _0057_ : _0060_;
  assign _0061_ = _T_4747 ? (* src = "crypto_accelerator.v:6346" *) io_dataIn[79:72] : matrix_1_2;
  assign _0062_ = _T_4775 ? (* src = "crypto_accelerator.v:6341" *) xorOut_1_2 : MixColsModule_io_out_1_2;
  assign _0063_ = state[0] ? (* src = "crypto_accelerator.v:6339" *) _0062_ : { _T_1963, _T_1964, _T_1965, _T_1966, _T_1967, _T_1968, _T_1969, _T_1970 };
  assign _0064_ = _T_4771 ? (* src = "crypto_accelerator.v:6337" *) _T_4726[79:72] : _0063_;
  assign _0007_ = io_ready ? (* src = "crypto_accelerator.v:6336" *) _0061_ : _0064_;
  assign _0065_ = _T_4747 ? (* src = "crypto_accelerator.v:6333" *) io_dataIn[87:80] : matrix_1_1;
  assign _0066_ = _T_4775 ? (* src = "crypto_accelerator.v:6328" *) xorOut_1_1 : MixColsModule_io_out_1_1;
  assign _0067_ = state[0] ? (* src = "crypto_accelerator.v:6326" *) _0066_ : { _T_1684, _T_1685, _T_1686, _T_1687, _T_1688, _T_1689, _T_1690, _T_1691 };
  assign _0068_ = _T_4771 ? (* src = "crypto_accelerator.v:6324" *) _T_4726[87:80] : _0067_;
  assign _0006_ = io_ready ? (* src = "crypto_accelerator.v:6323" *) _0065_ : _0068_;
  assign _0069_ = _T_4747 ? (* src = "crypto_accelerator.v:6320" *) io_dataIn[95:88] : matrix_1_0;
  assign _0070_ = _T_4775 ? (* src = "crypto_accelerator.v:6315" *) xorOut_1_0 : MixColsModule_io_out_1_0;
  assign _0071_ = state[0] ? (* src = "crypto_accelerator.v:6313" *) _0070_ : { _T_1405, _T_1406, _T_1407, _T_1408, _T_1409, _T_1410, _T_1411, _T_1412 };
  assign _0072_ = _T_4771 ? (* src = "crypto_accelerator.v:6311" *) _T_4726[95:88] : _0071_;
  assign _0005_ = io_ready ? (* src = "crypto_accelerator.v:6310" *) _0069_ : _0072_;
  assign _0073_ = _T_4747 ? (* src = "crypto_accelerator.v:6307" *) io_dataIn[103:96] : matrix_0_3;
  assign _0074_ = _T_4775 ? (* src = "crypto_accelerator.v:6302" *) xorOut_0_3 : MixColsModule_io_out_0_3;
  assign _0075_ = state[0] ? (* src = "crypto_accelerator.v:6300" *) _0074_ : { _T_1125, _T_1126, _T_1127, _T_1128, _T_1129, _T_1130, _T_1131, _T_1132 };
  assign _0076_ = _T_4771 ? (* src = "crypto_accelerator.v:6298" *) _T_4726[103:96] : _0075_;
  assign _0004_ = io_ready ? (* src = "crypto_accelerator.v:6297" *) _0073_ : _0076_;
  assign _0077_ = _T_4747 ? (* src = "crypto_accelerator.v:6294" *) io_dataIn[111:104] : matrix_0_2;
  assign _0078_ = _T_4775 ? (* src = "crypto_accelerator.v:6289" *) xorOut_0_2 : MixColsModule_io_out_0_2;
  assign _0079_ = state[0] ? (* src = "crypto_accelerator.v:6287" *) _0078_ : { _T_846, _T_847, _T_848, _T_849, _T_850, _T_851, _T_852, _T_853 };
  assign _0080_ = _T_4771 ? (* src = "crypto_accelerator.v:6285" *) _T_4726[111:104] : _0079_;
  assign _0003_ = io_ready ? (* src = "crypto_accelerator.v:6284" *) _0077_ : _0080_;
  assign _0081_ = _T_4747 ? (* src = "crypto_accelerator.v:6281" *) io_dataIn[119:112] : matrix_0_1;
  assign _0082_ = _T_4775 ? (* src = "crypto_accelerator.v:6276" *) xorOut_0_1 : MixColsModule_io_out_0_1;
  assign _0083_ = state[0] ? (* src = "crypto_accelerator.v:6274" *) _0082_ : { _T_567, _T_568, _T_569, _T_570, _T_571, _T_572, _T_573, _T_574 };
  assign _0084_ = _T_4771 ? (* src = "crypto_accelerator.v:6272" *) _T_4726[119:112] : _0083_;
  assign _0002_ = io_ready ? (* src = "crypto_accelerator.v:6271" *) _0081_ : _0084_;
  assign _0085_ = _T_4747 ? (* src = "crypto_accelerator.v:6268" *) io_dataIn[127:120] : matrix_0_0;
  assign _0086_ = _T_4775 ? (* src = "crypto_accelerator.v:6263" *) xorOut_0_0 : MixColsModule_io_out_0_0;
  assign _0087_ = state[0] ? (* src = "crypto_accelerator.v:6261" *) _0086_ : { _T_288, _T_289, _T_290, _T_291, _T_292, _T_293, _T_294, _T_295 };
  assign _0088_ = _T_4771 ? (* src = "crypto_accelerator.v:6259" *) _T_4726[127:120] : _0087_;
  assign _0001_ = io_ready ? (* src = "crypto_accelerator.v:6258" *) _0085_ : _0088_;
  assign _0089_ = _T_4747 ? (* src = "crypto_accelerator.v:6252" *) { 2'b01, _GEN_327 } : state;
  assign _0090_ = io_ready ? (* src = "crypto_accelerator.v:6250" *) _0089_ : _T_4778;
  assign _0017_ = reset ? (* src = "crypto_accelerator.v:6248" *) 6'b011110 : _0090_;
  assign _T_4778 = state - (* src = "crypto_accelerator.v:6111" *) 1'b1;
  assign keyEndAddr = io_aes256 ? (* src = "crypto_accelerator.v:5706" *) 3'b110 : 3'b010;
  assign _GEN_128 = _0018_ ? (* src = "crypto_accelerator.v:5819" *) io_keys_8_0_0 : io_keys_0_0_0;
  assign _GEN_129 = _0018_ ? (* src = "crypto_accelerator.v:5820" *) io_keys_8_0_1 : io_keys_0_0_1;
  assign _GEN_130 = _0018_ ? (* src = "crypto_accelerator.v:5821" *) io_keys_8_0_2 : io_keys_0_0_2;
  assign _GEN_131 = _0018_ ? (* src = "crypto_accelerator.v:5822" *) io_keys_8_0_3 : io_keys_0_0_3;
  assign _GEN_132 = _0018_ ? (* src = "crypto_accelerator.v:5823" *) io_keys_8_1_0 : io_keys_0_1_0;
  assign _GEN_133 = _0018_ ? (* src = "crypto_accelerator.v:5824" *) io_keys_8_1_1 : io_keys_0_1_1;
  assign _GEN_134 = _0018_ ? (* src = "crypto_accelerator.v:5825" *) io_keys_8_1_2 : io_keys_0_1_2;
  assign _GEN_135 = _0018_ ? (* src = "crypto_accelerator.v:5826" *) io_keys_8_1_3 : io_keys_0_1_3;
  assign _GEN_136 = _0018_ ? (* src = "crypto_accelerator.v:5827" *) io_keys_8_2_0 : io_keys_0_2_0;
  assign _GEN_137 = _0018_ ? (* src = "crypto_accelerator.v:5828" *) io_keys_8_2_1 : io_keys_0_2_1;
  assign _GEN_138 = _0018_ ? (* src = "crypto_accelerator.v:5829" *) io_keys_8_2_2 : io_keys_0_2_2;
  assign _GEN_139 = _0018_ ? (* src = "crypto_accelerator.v:5830" *) io_keys_8_2_3 : io_keys_0_2_3;
  assign _GEN_140 = _0018_ ? (* src = "crypto_accelerator.v:5831" *) io_keys_8_3_0 : io_keys_0_3_0;
  assign _GEN_141 = _0018_ ? (* src = "crypto_accelerator.v:5832" *) io_keys_8_3_1 : io_keys_0_3_1;
  assign _GEN_142 = _0018_ ? (* src = "crypto_accelerator.v:5833" *) io_keys_8_3_2 : io_keys_0_3_2;
  assign _GEN_143 = _0018_ ? (* src = "crypto_accelerator.v:5834" *) io_keys_8_3_3 : io_keys_0_3_3;
  assign _GEN_144 = _0019_ ? (* src = "crypto_accelerator.v:5835" *) io_keys_9_0_0 : _GEN_128;
  assign _GEN_145 = _0019_ ? (* src = "crypto_accelerator.v:5836" *) io_keys_9_0_1 : _GEN_129;
  assign _GEN_146 = _0019_ ? (* src = "crypto_accelerator.v:5837" *) io_keys_9_0_2 : _GEN_130;
  assign _GEN_147 = _0019_ ? (* src = "crypto_accelerator.v:5838" *) io_keys_9_0_3 : _GEN_131;
  assign _GEN_148 = _0019_ ? (* src = "crypto_accelerator.v:5839" *) io_keys_9_1_0 : _GEN_132;
  assign _GEN_149 = _0019_ ? (* src = "crypto_accelerator.v:5840" *) io_keys_9_1_1 : _GEN_133;
  assign _GEN_150 = _0019_ ? (* src = "crypto_accelerator.v:5841" *) io_keys_9_1_2 : _GEN_134;
  assign _GEN_151 = _0019_ ? (* src = "crypto_accelerator.v:5842" *) io_keys_9_1_3 : _GEN_135;
  assign _GEN_152 = _0019_ ? (* src = "crypto_accelerator.v:5843" *) io_keys_9_2_0 : _GEN_136;
  assign _GEN_153 = _0019_ ? (* src = "crypto_accelerator.v:5844" *) io_keys_9_2_1 : _GEN_137;
  assign _GEN_154 = _0019_ ? (* src = "crypto_accelerator.v:5845" *) io_keys_9_2_2 : _GEN_138;
  assign _GEN_155 = _0019_ ? (* src = "crypto_accelerator.v:5846" *) io_keys_9_2_3 : _GEN_139;
  assign _GEN_156 = _0019_ ? (* src = "crypto_accelerator.v:5847" *) io_keys_9_3_0 : _GEN_140;
  assign _GEN_157 = _0019_ ? (* src = "crypto_accelerator.v:5848" *) io_keys_9_3_1 : _GEN_141;
  assign _GEN_158 = _0019_ ? (* src = "crypto_accelerator.v:5849" *) io_keys_9_3_2 : _GEN_142;
  assign _GEN_159 = _0019_ ? (* src = "crypto_accelerator.v:5850" *) io_keys_9_3_3 : _GEN_143;
  assign _GEN_160 = _0020_ ? (* src = "crypto_accelerator.v:5851" *) io_keys_10_0_0 : _GEN_144;
  assign _GEN_161 = _0020_ ? (* src = "crypto_accelerator.v:5852" *) io_keys_10_0_1 : _GEN_145;
  assign _GEN_162 = _0020_ ? (* src = "crypto_accelerator.v:5853" *) io_keys_10_0_2 : _GEN_146;
  assign _GEN_163 = _0020_ ? (* src = "crypto_accelerator.v:5854" *) io_keys_10_0_3 : _GEN_147;
  assign _GEN_164 = _0020_ ? (* src = "crypto_accelerator.v:5855" *) io_keys_10_1_0 : _GEN_148;
  assign _GEN_165 = _0020_ ? (* src = "crypto_accelerator.v:5856" *) io_keys_10_1_1 : _GEN_149;
  assign _GEN_166 = _0020_ ? (* src = "crypto_accelerator.v:5857" *) io_keys_10_1_2 : _GEN_150;
  assign _GEN_167 = _0020_ ? (* src = "crypto_accelerator.v:5858" *) io_keys_10_1_3 : _GEN_151;
  assign _GEN_168 = _0020_ ? (* src = "crypto_accelerator.v:5859" *) io_keys_10_2_0 : _GEN_152;
  assign _GEN_169 = _0020_ ? (* src = "crypto_accelerator.v:5860" *) io_keys_10_2_1 : _GEN_153;
  assign _GEN_170 = _0020_ ? (* src = "crypto_accelerator.v:5861" *) io_keys_10_2_2 : _GEN_154;
  assign _GEN_171 = _0020_ ? (* src = "crypto_accelerator.v:5862" *) io_keys_10_2_3 : _GEN_155;
  assign _GEN_172 = _0020_ ? (* src = "crypto_accelerator.v:5863" *) io_keys_10_3_0 : _GEN_156;
  assign _GEN_173 = _0020_ ? (* src = "crypto_accelerator.v:5864" *) io_keys_10_3_1 : _GEN_157;
  assign _GEN_174 = _0020_ ? (* src = "crypto_accelerator.v:5865" *) io_keys_10_3_2 : _GEN_158;
  assign _GEN_175 = _0020_ ? (* src = "crypto_accelerator.v:5866" *) io_keys_10_3_3 : _GEN_159;
  assign _GEN_176 = _0021_ ? (* src = "crypto_accelerator.v:5867" *) io_keys_11_0_0 : _GEN_160;
  assign _GEN_177 = _0021_ ? (* src = "crypto_accelerator.v:5868" *) io_keys_11_0_1 : _GEN_161;
  assign _GEN_178 = _0021_ ? (* src = "crypto_accelerator.v:5869" *) io_keys_11_0_2 : _GEN_162;
  assign _GEN_179 = _0021_ ? (* src = "crypto_accelerator.v:5870" *) io_keys_11_0_3 : _GEN_163;
  assign _GEN_180 = _0021_ ? (* src = "crypto_accelerator.v:5871" *) io_keys_11_1_0 : _GEN_164;
  assign _GEN_181 = _0021_ ? (* src = "crypto_accelerator.v:5872" *) io_keys_11_1_1 : _GEN_165;
  assign _GEN_182 = _0021_ ? (* src = "crypto_accelerator.v:5873" *) io_keys_11_1_2 : _GEN_166;
  assign _GEN_183 = _0021_ ? (* src = "crypto_accelerator.v:5874" *) io_keys_11_1_3 : _GEN_167;
  assign _GEN_184 = _0021_ ? (* src = "crypto_accelerator.v:5875" *) io_keys_11_2_0 : _GEN_168;
  assign _GEN_185 = _0021_ ? (* src = "crypto_accelerator.v:5876" *) io_keys_11_2_1 : _GEN_169;
  assign _GEN_186 = _0021_ ? (* src = "crypto_accelerator.v:5877" *) io_keys_11_2_2 : _GEN_170;
  assign _GEN_187 = _0021_ ? (* src = "crypto_accelerator.v:5878" *) io_keys_11_2_3 : _GEN_171;
  assign _GEN_188 = _0021_ ? (* src = "crypto_accelerator.v:5879" *) io_keys_11_3_0 : _GEN_172;
  assign _GEN_189 = _0021_ ? (* src = "crypto_accelerator.v:5880" *) io_keys_11_3_1 : _GEN_173;
  assign _GEN_190 = _0021_ ? (* src = "crypto_accelerator.v:5881" *) io_keys_11_3_2 : _GEN_174;
  assign _GEN_191 = _0021_ ? (* src = "crypto_accelerator.v:5882" *) io_keys_11_3_3 : _GEN_175;
  assign _GEN_192 = _0022_ ? (* src = "crypto_accelerator.v:5883" *) io_keys_12_0_0 : _GEN_176;
  assign _GEN_193 = _0022_ ? (* src = "crypto_accelerator.v:5884" *) io_keys_12_0_1 : _GEN_177;
  assign _GEN_194 = _0022_ ? (* src = "crypto_accelerator.v:5885" *) io_keys_12_0_2 : _GEN_178;
  assign _GEN_195 = _0022_ ? (* src = "crypto_accelerator.v:5886" *) io_keys_12_0_3 : _GEN_179;
  assign _GEN_196 = _0022_ ? (* src = "crypto_accelerator.v:5887" *) io_keys_12_1_0 : _GEN_180;
  assign _GEN_197 = _0022_ ? (* src = "crypto_accelerator.v:5888" *) io_keys_12_1_1 : _GEN_181;
  assign _GEN_198 = _0022_ ? (* src = "crypto_accelerator.v:5889" *) io_keys_12_1_2 : _GEN_182;
  assign _GEN_199 = _0022_ ? (* src = "crypto_accelerator.v:5890" *) io_keys_12_1_3 : _GEN_183;
  assign _GEN_200 = _0022_ ? (* src = "crypto_accelerator.v:5891" *) io_keys_12_2_0 : _GEN_184;
  assign _GEN_201 = _0022_ ? (* src = "crypto_accelerator.v:5892" *) io_keys_12_2_1 : _GEN_185;
  assign _GEN_202 = _0022_ ? (* src = "crypto_accelerator.v:5893" *) io_keys_12_2_2 : _GEN_186;
  assign _GEN_203 = _0022_ ? (* src = "crypto_accelerator.v:5894" *) io_keys_12_2_3 : _GEN_187;
  assign _GEN_204 = _0022_ ? (* src = "crypto_accelerator.v:5895" *) io_keys_12_3_0 : _GEN_188;
  assign _GEN_205 = _0022_ ? (* src = "crypto_accelerator.v:5896" *) io_keys_12_3_1 : _GEN_189;
  assign _GEN_206 = _0022_ ? (* src = "crypto_accelerator.v:5897" *) io_keys_12_3_2 : _GEN_190;
  assign _GEN_207 = _0022_ ? (* src = "crypto_accelerator.v:5898" *) io_keys_12_3_3 : _GEN_191;
  assign _GEN_208 = _0023_ ? (* src = "crypto_accelerator.v:5899" *) io_keys_13_0_0 : _GEN_192;
  assign _GEN_209 = _0023_ ? (* src = "crypto_accelerator.v:5900" *) io_keys_13_0_1 : _GEN_193;
  assign _GEN_210 = _0023_ ? (* src = "crypto_accelerator.v:5901" *) io_keys_13_0_2 : _GEN_194;
  assign _GEN_211 = _0023_ ? (* src = "crypto_accelerator.v:5902" *) io_keys_13_0_3 : _GEN_195;
  assign _GEN_212 = _0023_ ? (* src = "crypto_accelerator.v:5903" *) io_keys_13_1_0 : _GEN_196;
  assign _GEN_213 = _0023_ ? (* src = "crypto_accelerator.v:5904" *) io_keys_13_1_1 : _GEN_197;
  assign _GEN_214 = _0023_ ? (* src = "crypto_accelerator.v:5905" *) io_keys_13_1_2 : _GEN_198;
  assign _GEN_215 = _0023_ ? (* src = "crypto_accelerator.v:5906" *) io_keys_13_1_3 : _GEN_199;
  assign _GEN_216 = _0023_ ? (* src = "crypto_accelerator.v:5907" *) io_keys_13_2_0 : _GEN_200;
  assign _GEN_217 = _0023_ ? (* src = "crypto_accelerator.v:5908" *) io_keys_13_2_1 : _GEN_201;
  assign _GEN_218 = _0023_ ? (* src = "crypto_accelerator.v:5909" *) io_keys_13_2_2 : _GEN_202;
  assign _GEN_219 = _0023_ ? (* src = "crypto_accelerator.v:5910" *) io_keys_13_2_3 : _GEN_203;
  assign _GEN_220 = _0023_ ? (* src = "crypto_accelerator.v:5911" *) io_keys_13_3_0 : _GEN_204;
  assign _GEN_221 = _0023_ ? (* src = "crypto_accelerator.v:5912" *) io_keys_13_3_1 : _GEN_205;
  assign _GEN_222 = _0023_ ? (* src = "crypto_accelerator.v:5913" *) io_keys_13_3_2 : _GEN_206;
  assign _GEN_223 = _0023_ ? (* src = "crypto_accelerator.v:5914" *) io_keys_13_3_3 : _GEN_207;
  assign _GEN_224 = _0024_ ? (* src = "crypto_accelerator.v:5915" *) io_keys_14_0_0 : _GEN_208;
  assign _GEN_225 = _0024_ ? (* src = "crypto_accelerator.v:5916" *) io_keys_14_0_1 : _GEN_209;
  assign _GEN_226 = _0024_ ? (* src = "crypto_accelerator.v:5917" *) io_keys_14_0_2 : _GEN_210;
  assign _GEN_227 = _0024_ ? (* src = "crypto_accelerator.v:5918" *) io_keys_14_0_3 : _GEN_211;
  assign _GEN_228 = _0024_ ? (* src = "crypto_accelerator.v:5919" *) io_keys_14_1_0 : _GEN_212;
  assign _GEN_229 = _0024_ ? (* src = "crypto_accelerator.v:5920" *) io_keys_14_1_1 : _GEN_213;
  assign _GEN_230 = _0024_ ? (* src = "crypto_accelerator.v:5921" *) io_keys_14_1_2 : _GEN_214;
  assign _GEN_231 = _0024_ ? (* src = "crypto_accelerator.v:5922" *) io_keys_14_1_3 : _GEN_215;
  assign _GEN_232 = _0024_ ? (* src = "crypto_accelerator.v:5923" *) io_keys_14_2_0 : _GEN_216;
  assign _GEN_233 = _0024_ ? (* src = "crypto_accelerator.v:5924" *) io_keys_14_2_1 : _GEN_217;
  assign _GEN_234 = _0024_ ? (* src = "crypto_accelerator.v:5925" *) io_keys_14_2_2 : _GEN_218;
  assign _GEN_235 = _0024_ ? (* src = "crypto_accelerator.v:5926" *) io_keys_14_2_3 : _GEN_219;
  assign _GEN_236 = _0024_ ? (* src = "crypto_accelerator.v:5927" *) io_keys_14_3_0 : _GEN_220;
  assign _GEN_237 = _0024_ ? (* src = "crypto_accelerator.v:5928" *) io_keys_14_3_1 : _GEN_221;
  assign _GEN_238 = _0024_ ? (* src = "crypto_accelerator.v:5929" *) io_keys_14_3_2 : _GEN_222;
  assign _GEN_239 = _0024_ ? (* src = "crypto_accelerator.v:5930" *) io_keys_14_3_3 : _GEN_223;
  assign _T_4541 = _T_4536 ? (* src = "crypto_accelerator.v:5953" *) _T_4539 : { _T_4534, 1'b0 };
  assign _T_4548 = _T_4543 ? (* src = "crypto_accelerator.v:5959" *) _T_4546 : { _T_4541[6:0], 1'b0 };
  assign _T_4556 = _T_4551 ? (* src = "crypto_accelerator.v:5966" *) _T_4554 : { _T_4549, 1'b0 };
  assign _T_4563 = _T_4558 ? (* src = "crypto_accelerator.v:5972" *) _T_4561 : { _T_4556[6:0], 1'b0 };
  assign _T_4575 = _T_4570 ? (* src = "crypto_accelerator.v:5987" *) _T_4573 : { _T_4568, 1'b0 };
  assign _T_4582[7:0] = _T_4577 ? (* src = "crypto_accelerator.v:5993" *) _T_4580 : { _T_4575[6:0], 1'b0 };
  assign _T_4590 = _T_4585 ? (* src = "crypto_accelerator.v:6000" *) _T_4588 : { _T_4583, 1'b0 };
  assign _T_4597 = _T_4592 ? (* src = "crypto_accelerator.v:6006" *) _T_4595[7:0] : { _T_4590[6:0], 1'b0 };
  assign _T_4609 = _T_4604 ? (* src = "crypto_accelerator.v:6021" *) _T_4607 : { _T_4602, 1'b0 };
  assign _T_4616[7:0] = _T_4611 ? (* src = "crypto_accelerator.v:6027" *) _T_4614 : { _T_4609[6:0], 1'b0 };
  assign _T_4624 = _T_4619 ? (* src = "crypto_accelerator.v:6034" *) _T_4622 : { _T_4617, 1'b0 };
  assign _T_4631[7:0] = _T_4626 ? (* src = "crypto_accelerator.v:6040" *) _T_4629[7:0] : { _T_4624[6:0], 1'b0 };
  assign _T_4643 = _T_4638 ? (* src = "crypto_accelerator.v:6055" *) _T_4641 : { _T_4636, 1'b0 };
  assign _T_4650[7:0] = _T_4645 ? (* src = "crypto_accelerator.v:6061" *) _T_4648 : { _T_4643[6:0], 1'b0 };
  assign _T_4658 = _T_4653 ? (* src = "crypto_accelerator.v:6068" *) _T_4656 : { _T_4651, 1'b0 };
  assign _T_4665 = _T_4660 ? (* src = "crypto_accelerator.v:6074" *) _T_4663[7:0] : { _T_4658[6:0], 1'b0 };
  assign _GEN_327 = io_aes256 ? (* src = "crypto_accelerator.v:6103" *) 4'b1101 : 4'b0101;
  assign _T_41 = matrix_0_0[7] ^ (* src = "crypto_accelerator.v:3498" *) matrix_0_0[4];
  assign _T_43 = matrix_0_0[6] ^ (* src = "crypto_accelerator.v:3499" *) matrix_0_0[4];
  assign _T_46 = matrix_0_0[7] ^ (* src = "crypto_accelerator.v:3501" *) matrix_0_0[6];
  assign _T_49 = matrix_0_0[4] ^ (* src = "crypto_accelerator.v:3503" *) matrix_0_0[3];
  assign _T_51 = matrix_0_0[3] ^ (* src = "crypto_accelerator.v:3504" *) matrix_0_0[0];
  assign _T_54 = matrix_0_0[1] ^ (* src = "crypto_accelerator.v:3506" *) matrix_0_0[0];
  assign _T_56 = matrix_0_0[6] ^ (* src = "crypto_accelerator.v:3507" *) _T_41;
  assign _T_59 = _T_44 ^ (* src = "crypto_accelerator.v:3509" *) _T_54;
  assign _T_61 = matrix_0_0[0] ^ (* src = "crypto_accelerator.v:3510" *) _T_49;
  assign _T_64 = _T_47 ^ (* src = "crypto_accelerator.v:3512" *) _T_52;
  assign _T_66 = _T_47 ^ (* src = "crypto_accelerator.v:3513" *) _T_54;
  assign _T_68 = _T_49 ^ (* src = "crypto_accelerator.v:3514" *) _T_54;
  assign _T_70 = matrix_0_0[5] ^ (* src = "crypto_accelerator.v:3515" *) _T_49;
  assign _T_73 = matrix_0_0[6] ^ (* src = "crypto_accelerator.v:3517" *) matrix_0_0[1];
  assign _T_75 = matrix_0_0[5] ^ (* src = "crypto_accelerator.v:3518" *) _T_59;
  assign _T_78 = _T_52 ^ (* src = "crypto_accelerator.v:3520" *) _T_73;
  assign _T_80 = matrix_0_0[3] ^ (* src = "crypto_accelerator.v:3521" *) _T_57;
  assign _T_82 = matrix_0_0[5] ^ (* src = "crypto_accelerator.v:3522" *) matrix_0_0[2];
  assign _T_85 = matrix_0_0[2] ^ (* src = "crypto_accelerator.v:3524" *) matrix_0_0[1];
  assign _T_88 = matrix_0_0[5] ^ (* src = "crypto_accelerator.v:3526" *) matrix_0_0[3];
  assign _T_91 = matrix_0_0[7] ^ (* src = "crypto_accelerator.v:3528" *) _T_83;
  assign _T_93 = _T_44 ^ (* src = "crypto_accelerator.v:3529" *) _T_83;
  assign _T_95 = _T_73 ^ (* src = "crypto_accelerator.v:3530" *) _T_89;
  assign _T_97 = _T_49 ^ (* src = "crypto_accelerator.v:3531" *) _T_86;
  assign _T_99 = _T_64 ^ (* src = "crypto_accelerator.v:3532" *) _T_97;
  assign _T_101 = _T_64 ^ (* src = "crypto_accelerator.v:3533" *) _T_86;
  assign _T_103 = _T_68 ^ (* src = "crypto_accelerator.v:3534" *) _T_95;
  assign _T_109 = _T_101 ^ (* src = "crypto_accelerator.v:3537" *) _T_105;
  assign _T_113 = _T_111 ^ (* src = "crypto_accelerator.v:3539" *) _T_105;
  assign _T_119 = _T_103 ^ (* src = "crypto_accelerator.v:3542" *) _T_115;
  assign _T_123 = _T_121 ^ (* src = "crypto_accelerator.v:3544" *) _T_115;
  assign _T_129 = _T_127 ^ (* src = "crypto_accelerator.v:3547" *) _T_125;
  assign _T_133 = _T_131 ^ (* src = "crypto_accelerator.v:3549" *) _T_125;
  assign _T_135 = _T_109 ^ (* src = "crypto_accelerator.v:3550" *) _T_107;
  assign _T_137 = _T_113 ^ (* src = "crypto_accelerator.v:3551" *) _T_52;
  assign _T_139 = _T_119 ^ (* src = "crypto_accelerator.v:3552" *) _T_117;
  assign _T_141 = _T_123 ^ (* src = "crypto_accelerator.v:3553" *) _T_133;
  assign _T_143 = _T_135 ^ (* src = "crypto_accelerator.v:3554" *) _T_129;
  assign _T_145 = _T_137 ^ (* src = "crypto_accelerator.v:3555" *) _T_133;
  assign _T_147 = _T_139 ^ (* src = "crypto_accelerator.v:3556" *) _T_129;
  assign _T_149 = _T_141 ^ (* src = "crypto_accelerator.v:3557" *) _T_71;
  assign _T_151 = _T_147 ^ (* src = "crypto_accelerator.v:3558" *) _T_149;
  assign _T_155 = _T_145 ^ (* src = "crypto_accelerator.v:3560" *) _T_153;
  assign _T_157 = _T_143 ^ (* src = "crypto_accelerator.v:3561" *) _T_145;
  assign _T_159 = _T_149 ^ (* src = "crypto_accelerator.v:3562" *) _T_153;
  assign _T_169 = _T_157 ^ (* src = "crypto_accelerator.v:3567" *) _T_153;
  assign _T_175 = _T_151 ^ (* src = "crypto_accelerator.v:3570" *) _T_153;
  assign _T_177 = _T_145 ^ (* src = "crypto_accelerator.v:3571" *) _T_161;
  assign _T_179 = _T_167 ^ (* src = "crypto_accelerator.v:3572" *) _T_169;
  assign _T_181 = _T_149 ^ (* src = "crypto_accelerator.v:3573" *) _T_163;
  assign _T_183 = _T_173 ^ (* src = "crypto_accelerator.v:3574" *) _T_175;
  assign _T_185 = _T_179 ^ (* src = "crypto_accelerator.v:3575" *) _T_183;
  assign _T_187 = _T_177 ^ (* src = "crypto_accelerator.v:3576" *) _T_181;
  assign _T_189 = _T_177 ^ (* src = "crypto_accelerator.v:3577" *) _T_179;
  assign _T_191 = _T_181 ^ (* src = "crypto_accelerator.v:3578" *) _T_183;
  assign _T_193 = _T_187 ^ (* src = "crypto_accelerator.v:3579" *) _T_185;
  assign _T_231 = _T_207 ^ (* src = "crypto_accelerator.v:3598" *) _T_225;
  assign _T_233 = _T_219 ^ (* src = "crypto_accelerator.v:3599" *) _T_221;
  assign _T_235 = _T_211 ^ (* src = "crypto_accelerator.v:3600" *) _T_227;
  assign _T_237 = _T_197 ^ (* src = "crypto_accelerator.v:3601" *) _T_203;
  assign _T_239 = _T_199 ^ (* src = "crypto_accelerator.v:3602" *) _T_215;
  assign _T_241 = _T_195 ^ (* src = "crypto_accelerator.v:3603" *) _T_205;
  assign _T_243 = _T_201 ^ (* src = "crypto_accelerator.v:3604" *) _T_223;
  assign _T_245 = _T_231 ^ (* src = "crypto_accelerator.v:3605" *) _T_233;
  assign _T_247 = _T_203 ^ (* src = "crypto_accelerator.v:3606" *) _T_209;
  assign _T_249 = _T_213 ^ (* src = "crypto_accelerator.v:3607" *) _T_229;
  assign _T_251 = _T_217 ^ (* src = "crypto_accelerator.v:3608" *) _T_239;
  assign _T_253 = _T_231 ^ (* src = "crypto_accelerator.v:3609" *) _T_237;
  assign _T_255 = _T_195 ^ (* src = "crypto_accelerator.v:3610" *) _T_199;
  assign _T_257 = _T_201 ^ (* src = "crypto_accelerator.v:3611" *) _T_205;
  assign _T_259 = _T_201 ^ (* src = "crypto_accelerator.v:3612" *) _T_227;
  assign _T_261 = _T_211 ^ (* src = "crypto_accelerator.v:3613" *) _T_221;
  assign _T_263 = _T_217 ^ (* src = "crypto_accelerator.v:3614" *) _T_225;
  assign _T_265 = _T_219 ^ (* src = "crypto_accelerator.v:3615" *) _T_235;
  assign _T_267 = _T_229 ^ (* src = "crypto_accelerator.v:3616" *) _T_241;
  assign _T_269 = _T_235 ^ (* src = "crypto_accelerator.v:3617" *) _T_237;
  assign _T_271 = _T_239 ^ (* src = "crypto_accelerator.v:3618" *) _T_243;
  assign _T_273 = _T_235 ^ (* src = "crypto_accelerator.v:3619" *) _T_245;
  assign _T_275 = _T_245 ^ (* src = "crypto_accelerator.v:3620" *) _T_247;
  assign _T_277 = _T_241 ^ (* src = "crypto_accelerator.v:3621" *) _T_245;
  assign _T_279 = _T_243 ^ (* src = "crypto_accelerator.v:3622" *) _T_251;
  assign _T_281 = _T_249 ^ (* src = "crypto_accelerator.v:3623" *) _T_253;
  assign _T_283 = _T_251 ^ (* src = "crypto_accelerator.v:3624" *) _T_267;
  assign _T_285 = _T_253 ^ (* src = "crypto_accelerator.v:3625" *) _T_279;
  assign _T_287 = _T_261 ^ (* src = "crypto_accelerator.v:3626" *) _T_271;
  assign _T_288 = _T_257 ^ (* src = "crypto_accelerator.v:3627" *) _T_273;
  assign _T_289 = _T_281 ^ (* src = "crypto_accelerator.v:3628" *) _T_287;
  assign _T_290 = _T_265 ^ (* src = "crypto_accelerator.v:3629" *) _T_285;
  assign _T_291 = _T_255 ^ (* src = "crypto_accelerator.v:3630" *) _T_273;
  assign _T_292 = _T_275 ^ (* src = "crypto_accelerator.v:3631" *) _T_283;
  assign _T_293 = _T_269 ^ (* src = "crypto_accelerator.v:3632" *) _T_277;
  assign _T_294 = _T_259 ^ (* src = "crypto_accelerator.v:3633" *) _T_275;
  assign _T_295 = _T_249 ^ (* src = "crypto_accelerator.v:3634" *) _T_263;
  assign _T_320 = matrix_3_1[7] ^ (* src = "crypto_accelerator.v:3636" *) matrix_3_1[4];
  assign _T_322 = matrix_3_1[6] ^ (* src = "crypto_accelerator.v:3637" *) matrix_3_1[4];
  assign _T_325 = matrix_3_1[7] ^ (* src = "crypto_accelerator.v:3639" *) matrix_3_1[6];
  assign _T_328 = matrix_3_1[4] ^ (* src = "crypto_accelerator.v:3641" *) matrix_3_1[3];
  assign _T_330 = matrix_3_1[3] ^ (* src = "crypto_accelerator.v:3642" *) matrix_3_1[0];
  assign _T_333 = matrix_3_1[1] ^ (* src = "crypto_accelerator.v:3644" *) matrix_3_1[0];
  assign _T_335 = matrix_3_1[6] ^ (* src = "crypto_accelerator.v:3645" *) _T_320;
  assign _T_338 = _T_323 ^ (* src = "crypto_accelerator.v:3647" *) _T_333;
  assign _T_340 = matrix_3_1[0] ^ (* src = "crypto_accelerator.v:3648" *) _T_328;
  assign _T_343 = _T_326 ^ (* src = "crypto_accelerator.v:3650" *) _T_331;
  assign _T_345 = _T_326 ^ (* src = "crypto_accelerator.v:3651" *) _T_333;
  assign _T_347 = _T_328 ^ (* src = "crypto_accelerator.v:3652" *) _T_333;
  assign _T_349 = matrix_3_1[5] ^ (* src = "crypto_accelerator.v:3653" *) _T_328;
  assign _T_352 = matrix_3_1[6] ^ (* src = "crypto_accelerator.v:3655" *) matrix_3_1[1];
  assign _T_354 = matrix_3_1[5] ^ (* src = "crypto_accelerator.v:3656" *) _T_338;
  assign _T_357 = _T_331 ^ (* src = "crypto_accelerator.v:3658" *) _T_352;
  assign _T_359 = matrix_3_1[3] ^ (* src = "crypto_accelerator.v:3659" *) _T_336;
  assign _T_361 = matrix_3_1[5] ^ (* src = "crypto_accelerator.v:3660" *) matrix_3_1[2];
  assign _T_364 = matrix_3_1[2] ^ (* src = "crypto_accelerator.v:3662" *) matrix_3_1[1];
  assign _T_367 = matrix_3_1[5] ^ (* src = "crypto_accelerator.v:3664" *) matrix_3_1[3];
  assign _T_370 = matrix_3_1[7] ^ (* src = "crypto_accelerator.v:3666" *) _T_362;
  assign _T_372 = _T_323 ^ (* src = "crypto_accelerator.v:3667" *) _T_362;
  assign _T_374 = _T_352 ^ (* src = "crypto_accelerator.v:3668" *) _T_368;
  assign _T_376 = _T_328 ^ (* src = "crypto_accelerator.v:3669" *) _T_365;
  assign _T_378 = _T_343 ^ (* src = "crypto_accelerator.v:3670" *) _T_376;
  assign _T_380 = _T_343 ^ (* src = "crypto_accelerator.v:3671" *) _T_365;
  assign _T_382 = _T_347 ^ (* src = "crypto_accelerator.v:3672" *) _T_374;
  assign _T_388 = _T_380 ^ (* src = "crypto_accelerator.v:3675" *) _T_384;
  assign _T_392 = _T_390 ^ (* src = "crypto_accelerator.v:3677" *) _T_384;
  assign _T_398 = _T_382 ^ (* src = "crypto_accelerator.v:3680" *) _T_394;
  assign _T_402 = _T_400 ^ (* src = "crypto_accelerator.v:3682" *) _T_394;
  assign _T_408 = _T_406 ^ (* src = "crypto_accelerator.v:3685" *) _T_404;
  assign _T_412 = _T_410 ^ (* src = "crypto_accelerator.v:3687" *) _T_404;
  assign _T_414 = _T_388 ^ (* src = "crypto_accelerator.v:3688" *) _T_386;
  assign _T_416 = _T_392 ^ (* src = "crypto_accelerator.v:3689" *) _T_331;
  assign _T_418 = _T_398 ^ (* src = "crypto_accelerator.v:3690" *) _T_396;
  assign _T_420 = _T_402 ^ (* src = "crypto_accelerator.v:3691" *) _T_412;
  assign _T_422 = _T_414 ^ (* src = "crypto_accelerator.v:3692" *) _T_408;
  assign _T_424 = _T_416 ^ (* src = "crypto_accelerator.v:3693" *) _T_412;
  assign _T_426 = _T_418 ^ (* src = "crypto_accelerator.v:3694" *) _T_408;
  assign _T_428 = _T_420 ^ (* src = "crypto_accelerator.v:3695" *) _T_350;
  assign _T_430 = _T_426 ^ (* src = "crypto_accelerator.v:3696" *) _T_428;
  assign _T_434 = _T_424 ^ (* src = "crypto_accelerator.v:3698" *) _T_432;
  assign _T_436 = _T_422 ^ (* src = "crypto_accelerator.v:3699" *) _T_424;
  assign _T_438 = _T_428 ^ (* src = "crypto_accelerator.v:3700" *) _T_432;
  assign _T_448 = _T_436 ^ (* src = "crypto_accelerator.v:3705" *) _T_432;
  assign _T_454 = _T_430 ^ (* src = "crypto_accelerator.v:3708" *) _T_432;
  assign _T_456 = _T_424 ^ (* src = "crypto_accelerator.v:3709" *) _T_440;
  assign _T_458 = _T_446 ^ (* src = "crypto_accelerator.v:3710" *) _T_448;
  assign _T_460 = _T_428 ^ (* src = "crypto_accelerator.v:3711" *) _T_442;
  assign _T_462 = _T_452 ^ (* src = "crypto_accelerator.v:3712" *) _T_454;
  assign _T_464 = _T_458 ^ (* src = "crypto_accelerator.v:3713" *) _T_462;
  assign _T_466 = _T_456 ^ (* src = "crypto_accelerator.v:3714" *) _T_460;
  assign _T_468 = _T_456 ^ (* src = "crypto_accelerator.v:3715" *) _T_458;
  assign _T_470 = _T_460 ^ (* src = "crypto_accelerator.v:3716" *) _T_462;
  assign _T_472 = _T_466 ^ (* src = "crypto_accelerator.v:3717" *) _T_464;
  assign _T_510 = _T_486 ^ (* src = "crypto_accelerator.v:3736" *) _T_504;
  assign _T_512 = _T_498 ^ (* src = "crypto_accelerator.v:3737" *) _T_500;
  assign _T_514 = _T_490 ^ (* src = "crypto_accelerator.v:3738" *) _T_506;
  assign _T_516 = _T_476 ^ (* src = "crypto_accelerator.v:3739" *) _T_482;
  assign _T_518 = _T_478 ^ (* src = "crypto_accelerator.v:3740" *) _T_494;
  assign _T_520 = _T_474 ^ (* src = "crypto_accelerator.v:3741" *) _T_484;
  assign _T_522 = _T_480 ^ (* src = "crypto_accelerator.v:3742" *) _T_502;
  assign _T_524 = _T_510 ^ (* src = "crypto_accelerator.v:3743" *) _T_512;
  assign _T_526 = _T_482 ^ (* src = "crypto_accelerator.v:3744" *) _T_488;
  assign _T_528 = _T_492 ^ (* src = "crypto_accelerator.v:3745" *) _T_508;
  assign _T_530 = _T_496 ^ (* src = "crypto_accelerator.v:3746" *) _T_518;
  assign _T_532 = _T_510 ^ (* src = "crypto_accelerator.v:3747" *) _T_516;
  assign _T_534 = _T_474 ^ (* src = "crypto_accelerator.v:3748" *) _T_478;
  assign _T_536 = _T_480 ^ (* src = "crypto_accelerator.v:3749" *) _T_484;
  assign _T_538 = _T_480 ^ (* src = "crypto_accelerator.v:3750" *) _T_506;
  assign _T_540 = _T_490 ^ (* src = "crypto_accelerator.v:3751" *) _T_500;
  assign _T_542 = _T_496 ^ (* src = "crypto_accelerator.v:3752" *) _T_504;
  assign _T_544 = _T_498 ^ (* src = "crypto_accelerator.v:3753" *) _T_514;
  assign _T_546 = _T_508 ^ (* src = "crypto_accelerator.v:3754" *) _T_520;
  assign _T_548 = _T_514 ^ (* src = "crypto_accelerator.v:3755" *) _T_516;
  assign _T_550 = _T_518 ^ (* src = "crypto_accelerator.v:3756" *) _T_522;
  assign _T_552 = _T_514 ^ (* src = "crypto_accelerator.v:3757" *) _T_524;
  assign _T_554 = _T_524 ^ (* src = "crypto_accelerator.v:3758" *) _T_526;
  assign _T_556 = _T_520 ^ (* src = "crypto_accelerator.v:3759" *) _T_524;
  assign _T_558 = _T_522 ^ (* src = "crypto_accelerator.v:3760" *) _T_530;
  assign _T_560 = _T_528 ^ (* src = "crypto_accelerator.v:3761" *) _T_532;
  assign _T_562 = _T_530 ^ (* src = "crypto_accelerator.v:3762" *) _T_546;
  assign _T_564 = _T_532 ^ (* src = "crypto_accelerator.v:3763" *) _T_558;
  assign _T_566 = _T_540 ^ (* src = "crypto_accelerator.v:3764" *) _T_550;
  assign _T_567 = _T_536 ^ (* src = "crypto_accelerator.v:3765" *) _T_552;
  assign _T_568 = _T_560 ^ (* src = "crypto_accelerator.v:3766" *) _T_566;
  assign _T_569 = _T_544 ^ (* src = "crypto_accelerator.v:3767" *) _T_564;
  assign _T_570 = _T_534 ^ (* src = "crypto_accelerator.v:3768" *) _T_552;
  assign _T_571 = _T_554 ^ (* src = "crypto_accelerator.v:3769" *) _T_562;
  assign _T_572 = _T_548 ^ (* src = "crypto_accelerator.v:3770" *) _T_556;
  assign _T_573 = _T_538 ^ (* src = "crypto_accelerator.v:3771" *) _T_554;
  assign _T_574 = _T_528 ^ (* src = "crypto_accelerator.v:3772" *) _T_542;
  assign _T_599 = matrix_2_2[7] ^ (* src = "crypto_accelerator.v:3774" *) matrix_2_2[4];
  assign _T_601 = matrix_2_2[6] ^ (* src = "crypto_accelerator.v:3775" *) matrix_2_2[4];
  assign _T_604 = matrix_2_2[7] ^ (* src = "crypto_accelerator.v:3777" *) matrix_2_2[6];
  assign _T_607 = matrix_2_2[4] ^ (* src = "crypto_accelerator.v:3779" *) matrix_2_2[3];
  assign _T_609 = matrix_2_2[3] ^ (* src = "crypto_accelerator.v:3780" *) matrix_2_2[0];
  assign _T_612 = matrix_2_2[1] ^ (* src = "crypto_accelerator.v:3782" *) matrix_2_2[0];
  assign _T_614 = matrix_2_2[6] ^ (* src = "crypto_accelerator.v:3783" *) _T_599;
  assign _T_617 = _T_602 ^ (* src = "crypto_accelerator.v:3785" *) _T_612;
  assign _T_619 = matrix_2_2[0] ^ (* src = "crypto_accelerator.v:3786" *) _T_607;
  assign _T_622 = _T_605 ^ (* src = "crypto_accelerator.v:3788" *) _T_610;
  assign _T_624 = _T_605 ^ (* src = "crypto_accelerator.v:3789" *) _T_612;
  assign _T_626 = _T_607 ^ (* src = "crypto_accelerator.v:3790" *) _T_612;
  assign _T_628 = matrix_2_2[5] ^ (* src = "crypto_accelerator.v:3791" *) _T_607;
  assign _T_631 = matrix_2_2[6] ^ (* src = "crypto_accelerator.v:3793" *) matrix_2_2[1];
  assign _T_633 = matrix_2_2[5] ^ (* src = "crypto_accelerator.v:3794" *) _T_617;
  assign _T_636 = _T_610 ^ (* src = "crypto_accelerator.v:3796" *) _T_631;
  assign _T_638 = matrix_2_2[3] ^ (* src = "crypto_accelerator.v:3797" *) _T_615;
  assign _T_640 = matrix_2_2[5] ^ (* src = "crypto_accelerator.v:3798" *) matrix_2_2[2];
  assign _T_643 = matrix_2_2[2] ^ (* src = "crypto_accelerator.v:3800" *) matrix_2_2[1];
  assign _T_646 = matrix_2_2[5] ^ (* src = "crypto_accelerator.v:3802" *) matrix_2_2[3];
  assign _T_649 = matrix_2_2[7] ^ (* src = "crypto_accelerator.v:3804" *) _T_641;
  assign _T_651 = _T_602 ^ (* src = "crypto_accelerator.v:3805" *) _T_641;
  assign _T_653 = _T_631 ^ (* src = "crypto_accelerator.v:3806" *) _T_647;
  assign _T_655 = _T_607 ^ (* src = "crypto_accelerator.v:3807" *) _T_644;
  assign _T_657 = _T_622 ^ (* src = "crypto_accelerator.v:3808" *) _T_655;
  assign _T_659 = _T_622 ^ (* src = "crypto_accelerator.v:3809" *) _T_644;
  assign _T_661 = _T_626 ^ (* src = "crypto_accelerator.v:3810" *) _T_653;
  assign _T_667 = _T_659 ^ (* src = "crypto_accelerator.v:3813" *) _T_663;
  assign _T_671 = _T_669 ^ (* src = "crypto_accelerator.v:3815" *) _T_663;
  assign _T_677 = _T_661 ^ (* src = "crypto_accelerator.v:3818" *) _T_673;
  assign _T_681 = _T_679 ^ (* src = "crypto_accelerator.v:3820" *) _T_673;
  assign _T_687 = _T_685 ^ (* src = "crypto_accelerator.v:3823" *) _T_683;
  assign _T_691 = _T_689 ^ (* src = "crypto_accelerator.v:3825" *) _T_683;
  assign _T_693 = _T_667 ^ (* src = "crypto_accelerator.v:3826" *) _T_665;
  assign _T_695 = _T_671 ^ (* src = "crypto_accelerator.v:3827" *) _T_610;
  assign _T_697 = _T_677 ^ (* src = "crypto_accelerator.v:3828" *) _T_675;
  assign _T_699 = _T_681 ^ (* src = "crypto_accelerator.v:3829" *) _T_691;
  assign _T_701 = _T_693 ^ (* src = "crypto_accelerator.v:3830" *) _T_687;
  assign _T_703 = _T_695 ^ (* src = "crypto_accelerator.v:3831" *) _T_691;
  assign _T_705 = _T_697 ^ (* src = "crypto_accelerator.v:3832" *) _T_687;
  assign _T_707 = _T_699 ^ (* src = "crypto_accelerator.v:3833" *) _T_629;
  assign _T_709 = _T_705 ^ (* src = "crypto_accelerator.v:3834" *) _T_707;
  assign _T_713 = _T_703 ^ (* src = "crypto_accelerator.v:3836" *) _T_711;
  assign _T_715 = _T_701 ^ (* src = "crypto_accelerator.v:3837" *) _T_703;
  assign _T_717 = _T_707 ^ (* src = "crypto_accelerator.v:3838" *) _T_711;
  assign _T_727 = _T_715 ^ (* src = "crypto_accelerator.v:3843" *) _T_711;
  assign _T_733 = _T_709 ^ (* src = "crypto_accelerator.v:3846" *) _T_711;
  assign _T_735 = _T_703 ^ (* src = "crypto_accelerator.v:3847" *) _T_719;
  assign _T_737 = _T_725 ^ (* src = "crypto_accelerator.v:3848" *) _T_727;
  assign _T_739 = _T_707 ^ (* src = "crypto_accelerator.v:3849" *) _T_721;
  assign _T_741 = _T_731 ^ (* src = "crypto_accelerator.v:3850" *) _T_733;
  assign _T_743 = _T_737 ^ (* src = "crypto_accelerator.v:3851" *) _T_741;
  assign _T_745 = _T_735 ^ (* src = "crypto_accelerator.v:3852" *) _T_739;
  assign _T_747 = _T_735 ^ (* src = "crypto_accelerator.v:3853" *) _T_737;
  assign _T_749 = _T_739 ^ (* src = "crypto_accelerator.v:3854" *) _T_741;
  assign _T_751 = _T_745 ^ (* src = "crypto_accelerator.v:3855" *) _T_743;
  assign _T_789 = _T_765 ^ (* src = "crypto_accelerator.v:3874" *) _T_783;
  assign _T_791 = _T_777 ^ (* src = "crypto_accelerator.v:3875" *) _T_779;
  assign _T_793 = _T_769 ^ (* src = "crypto_accelerator.v:3876" *) _T_785;
  assign _T_795 = _T_755 ^ (* src = "crypto_accelerator.v:3877" *) _T_761;
  assign _T_797 = _T_757 ^ (* src = "crypto_accelerator.v:3878" *) _T_773;
  assign _T_799 = _T_753 ^ (* src = "crypto_accelerator.v:3879" *) _T_763;
  assign _T_801 = _T_759 ^ (* src = "crypto_accelerator.v:3880" *) _T_781;
  assign _T_803 = _T_789 ^ (* src = "crypto_accelerator.v:3881" *) _T_791;
  assign _T_805 = _T_761 ^ (* src = "crypto_accelerator.v:3882" *) _T_767;
  assign _T_807 = _T_771 ^ (* src = "crypto_accelerator.v:3883" *) _T_787;
  assign _T_809 = _T_775 ^ (* src = "crypto_accelerator.v:3884" *) _T_797;
  assign _T_811 = _T_789 ^ (* src = "crypto_accelerator.v:3885" *) _T_795;
  assign _T_813 = _T_753 ^ (* src = "crypto_accelerator.v:3886" *) _T_757;
  assign _T_815 = _T_759 ^ (* src = "crypto_accelerator.v:3887" *) _T_763;
  assign _T_817 = _T_759 ^ (* src = "crypto_accelerator.v:3888" *) _T_785;
  assign _T_819 = _T_769 ^ (* src = "crypto_accelerator.v:3889" *) _T_779;
  assign _T_821 = _T_775 ^ (* src = "crypto_accelerator.v:3890" *) _T_783;
  assign _T_823 = _T_777 ^ (* src = "crypto_accelerator.v:3891" *) _T_793;
  assign _T_825 = _T_787 ^ (* src = "crypto_accelerator.v:3892" *) _T_799;
  assign _T_827 = _T_793 ^ (* src = "crypto_accelerator.v:3893" *) _T_795;
  assign _T_829 = _T_797 ^ (* src = "crypto_accelerator.v:3894" *) _T_801;
  assign _T_831 = _T_793 ^ (* src = "crypto_accelerator.v:3895" *) _T_803;
  assign _T_833 = _T_803 ^ (* src = "crypto_accelerator.v:3896" *) _T_805;
  assign _T_835 = _T_799 ^ (* src = "crypto_accelerator.v:3897" *) _T_803;
  assign _T_837 = _T_801 ^ (* src = "crypto_accelerator.v:3898" *) _T_809;
  assign _T_839 = _T_807 ^ (* src = "crypto_accelerator.v:3899" *) _T_811;
  assign _T_841 = _T_809 ^ (* src = "crypto_accelerator.v:3900" *) _T_825;
  assign _T_843 = _T_811 ^ (* src = "crypto_accelerator.v:3901" *) _T_837;
  assign _T_845 = _T_819 ^ (* src = "crypto_accelerator.v:3902" *) _T_829;
  assign _T_846 = _T_815 ^ (* src = "crypto_accelerator.v:3903" *) _T_831;
  assign _T_847 = _T_839 ^ (* src = "crypto_accelerator.v:3904" *) _T_845;
  assign _T_848 = _T_823 ^ (* src = "crypto_accelerator.v:3905" *) _T_843;
  assign _T_849 = _T_813 ^ (* src = "crypto_accelerator.v:3906" *) _T_831;
  assign _T_850 = _T_833 ^ (* src = "crypto_accelerator.v:3907" *) _T_841;
  assign _T_851 = _T_827 ^ (* src = "crypto_accelerator.v:3908" *) _T_835;
  assign _T_852 = _T_817 ^ (* src = "crypto_accelerator.v:3909" *) _T_833;
  assign _T_853 = _T_807 ^ (* src = "crypto_accelerator.v:3910" *) _T_821;
  assign _T_878 = matrix_1_3[7] ^ (* src = "crypto_accelerator.v:3912" *) matrix_1_3[4];
  assign _T_880 = matrix_1_3[6] ^ (* src = "crypto_accelerator.v:3913" *) matrix_1_3[4];
  assign _T_883 = matrix_1_3[7] ^ (* src = "crypto_accelerator.v:3915" *) matrix_1_3[6];
  assign _T_886 = matrix_1_3[4] ^ (* src = "crypto_accelerator.v:3917" *) matrix_1_3[3];
  assign _T_888 = matrix_1_3[3] ^ (* src = "crypto_accelerator.v:3918" *) matrix_1_3[0];
  assign _T_891 = matrix_1_3[1] ^ (* src = "crypto_accelerator.v:3920" *) matrix_1_3[0];
  assign _T_893 = matrix_1_3[6] ^ (* src = "crypto_accelerator.v:3921" *) _T_878;
  assign _T_896 = _T_881 ^ (* src = "crypto_accelerator.v:3923" *) _T_891;
  assign _T_898 = matrix_1_3[0] ^ (* src = "crypto_accelerator.v:3924" *) _T_886;
  assign _T_901 = _T_884 ^ (* src = "crypto_accelerator.v:3926" *) _T_889;
  assign _T_903 = _T_884 ^ (* src = "crypto_accelerator.v:3927" *) _T_891;
  assign _T_905 = _T_886 ^ (* src = "crypto_accelerator.v:3928" *) _T_891;
  assign _T_907 = matrix_1_3[5] ^ (* src = "crypto_accelerator.v:3929" *) _T_886;
  assign _T_910 = matrix_1_3[6] ^ (* src = "crypto_accelerator.v:3931" *) matrix_1_3[1];
  assign _T_912 = matrix_1_3[5] ^ (* src = "crypto_accelerator.v:3932" *) _T_896;
  assign _T_915 = _T_889 ^ (* src = "crypto_accelerator.v:3934" *) _T_910;
  assign _T_917 = matrix_1_3[3] ^ (* src = "crypto_accelerator.v:3935" *) _T_894;
  assign _T_919 = matrix_1_3[5] ^ (* src = "crypto_accelerator.v:3936" *) matrix_1_3[2];
  assign _T_922 = matrix_1_3[2] ^ (* src = "crypto_accelerator.v:3938" *) matrix_1_3[1];
  assign _T_925 = matrix_1_3[5] ^ (* src = "crypto_accelerator.v:3940" *) matrix_1_3[3];
  assign _T_928 = matrix_1_3[7] ^ (* src = "crypto_accelerator.v:3942" *) _T_920;
  assign _T_930 = _T_881 ^ (* src = "crypto_accelerator.v:3943" *) _T_920;
  assign _T_932 = _T_910 ^ (* src = "crypto_accelerator.v:3944" *) _T_926;
  assign _T_934 = _T_886 ^ (* src = "crypto_accelerator.v:3945" *) _T_923;
  assign _T_936 = _T_901 ^ (* src = "crypto_accelerator.v:3946" *) _T_934;
  assign _T_938 = _T_901 ^ (* src = "crypto_accelerator.v:3947" *) _T_923;
  assign _T_940 = _T_905 ^ (* src = "crypto_accelerator.v:3948" *) _T_932;
  assign _T_946 = _T_938 ^ (* src = "crypto_accelerator.v:3951" *) _T_942;
  assign _T_950 = _T_948 ^ (* src = "crypto_accelerator.v:3953" *) _T_942;
  assign _T_956 = _T_940 ^ (* src = "crypto_accelerator.v:3956" *) _T_952;
  assign _T_960 = _T_958 ^ (* src = "crypto_accelerator.v:3958" *) _T_952;
  assign _T_966 = _T_964 ^ (* src = "crypto_accelerator.v:3961" *) _T_962;
  assign _T_970 = _T_968 ^ (* src = "crypto_accelerator.v:3963" *) _T_962;
  assign _T_972 = _T_946 ^ (* src = "crypto_accelerator.v:3964" *) _T_944;
  assign _T_974 = _T_950 ^ (* src = "crypto_accelerator.v:3965" *) _T_889;
  assign _T_976 = _T_956 ^ (* src = "crypto_accelerator.v:3966" *) _T_954;
  assign _T_978 = _T_960 ^ (* src = "crypto_accelerator.v:3967" *) _T_970;
  assign _T_980 = _T_972 ^ (* src = "crypto_accelerator.v:3968" *) _T_966;
  assign _T_982 = _T_974 ^ (* src = "crypto_accelerator.v:3969" *) _T_970;
  assign _T_984 = _T_976 ^ (* src = "crypto_accelerator.v:3970" *) _T_966;
  assign _T_986 = _T_978 ^ (* src = "crypto_accelerator.v:3971" *) _T_908;
  assign _T_988 = _T_984 ^ (* src = "crypto_accelerator.v:3972" *) _T_986;
  assign _T_992 = _T_982 ^ (* src = "crypto_accelerator.v:3974" *) _T_990;
  assign _T_994 = _T_980 ^ (* src = "crypto_accelerator.v:3975" *) _T_982;
  assign _T_996 = _T_986 ^ (* src = "crypto_accelerator.v:3976" *) _T_990;
  assign _T_1006 = _T_994 ^ (* src = "crypto_accelerator.v:3981" *) _T_990;
  assign _T_1012 = _T_988 ^ (* src = "crypto_accelerator.v:3984" *) _T_990;
  assign _T_1014 = _T_982 ^ (* src = "crypto_accelerator.v:3985" *) _T_998;
  assign _T_1016 = _T_1004 ^ (* src = "crypto_accelerator.v:3986" *) _T_1006;
  assign _T_1018 = _T_986 ^ (* src = "crypto_accelerator.v:3987" *) _T_1000;
  assign _T_1020 = _T_1010 ^ (* src = "crypto_accelerator.v:3988" *) _T_1012;
  assign _T_1022 = _T_1016 ^ (* src = "crypto_accelerator.v:3989" *) _T_1020;
  assign _T_1024 = _T_1014 ^ (* src = "crypto_accelerator.v:3990" *) _T_1018;
  assign _T_1026 = _T_1014 ^ (* src = "crypto_accelerator.v:3991" *) _T_1016;
  assign _T_1028 = _T_1018 ^ (* src = "crypto_accelerator.v:3992" *) _T_1020;
  assign _T_1030 = _T_1024 ^ (* src = "crypto_accelerator.v:3993" *) _T_1022;
  assign _T_1068 = _T_1044 ^ (* src = "crypto_accelerator.v:4012" *) _T_1062;
  assign _T_1070 = _T_1056 ^ (* src = "crypto_accelerator.v:4013" *) _T_1058;
  assign _T_1072 = _T_1048 ^ (* src = "crypto_accelerator.v:4014" *) _T_1064;
  assign _T_1074 = _T_1034 ^ (* src = "crypto_accelerator.v:4015" *) _T_1040;
  assign _T_1076 = _T_1036 ^ (* src = "crypto_accelerator.v:4016" *) _T_1052;
  assign _T_1078 = _T_1032 ^ (* src = "crypto_accelerator.v:4017" *) _T_1042;
  assign _T_1080 = _T_1038 ^ (* src = "crypto_accelerator.v:4018" *) _T_1060;
  assign _T_1082 = _T_1068 ^ (* src = "crypto_accelerator.v:4019" *) _T_1070;
  assign _T_1084 = _T_1040 ^ (* src = "crypto_accelerator.v:4020" *) _T_1046;
  assign _T_1086 = _T_1050 ^ (* src = "crypto_accelerator.v:4021" *) _T_1066;
  assign _T_1088 = _T_1054 ^ (* src = "crypto_accelerator.v:4022" *) _T_1076;
  assign _T_1090 = _T_1068 ^ (* src = "crypto_accelerator.v:4023" *) _T_1074;
  assign _T_1092 = _T_1032 ^ (* src = "crypto_accelerator.v:4024" *) _T_1036;
  assign _T_1094 = _T_1038 ^ (* src = "crypto_accelerator.v:4025" *) _T_1042;
  assign _T_1096 = _T_1038 ^ (* src = "crypto_accelerator.v:4026" *) _T_1064;
  assign _T_1098 = _T_1048 ^ (* src = "crypto_accelerator.v:4027" *) _T_1058;
  assign _T_1100 = _T_1054 ^ (* src = "crypto_accelerator.v:4028" *) _T_1062;
  assign _T_1102 = _T_1056 ^ (* src = "crypto_accelerator.v:4029" *) _T_1072;
  assign _T_1104 = _T_1066 ^ (* src = "crypto_accelerator.v:4030" *) _T_1078;
  assign _T_1106 = _T_1072 ^ (* src = "crypto_accelerator.v:4031" *) _T_1074;
  assign _T_1108 = _T_1076 ^ (* src = "crypto_accelerator.v:4032" *) _T_1080;
  assign _T_1110 = _T_1072 ^ (* src = "crypto_accelerator.v:4033" *) _T_1082;
  assign _T_1112 = _T_1082 ^ (* src = "crypto_accelerator.v:4034" *) _T_1084;
  assign _T_1114 = _T_1078 ^ (* src = "crypto_accelerator.v:4035" *) _T_1082;
  assign _T_1116 = _T_1080 ^ (* src = "crypto_accelerator.v:4036" *) _T_1088;
  assign _T_1118 = _T_1086 ^ (* src = "crypto_accelerator.v:4037" *) _T_1090;
  assign _T_1120 = _T_1088 ^ (* src = "crypto_accelerator.v:4038" *) _T_1104;
  assign _T_1122 = _T_1090 ^ (* src = "crypto_accelerator.v:4039" *) _T_1116;
  assign _T_1124 = _T_1098 ^ (* src = "crypto_accelerator.v:4040" *) _T_1108;
  assign _T_1125 = _T_1094 ^ (* src = "crypto_accelerator.v:4041" *) _T_1110;
  assign _T_1126 = _T_1118 ^ (* src = "crypto_accelerator.v:4042" *) _T_1124;
  assign _T_1127 = _T_1102 ^ (* src = "crypto_accelerator.v:4043" *) _T_1122;
  assign _T_1128 = _T_1092 ^ (* src = "crypto_accelerator.v:4044" *) _T_1110;
  assign _T_1129 = _T_1112 ^ (* src = "crypto_accelerator.v:4045" *) _T_1120;
  assign _T_1130 = _T_1106 ^ (* src = "crypto_accelerator.v:4046" *) _T_1114;
  assign _T_1131 = _T_1096 ^ (* src = "crypto_accelerator.v:4047" *) _T_1112;
  assign _T_1132 = _T_1086 ^ (* src = "crypto_accelerator.v:4048" *) _T_1100;
  assign _T_1158 = matrix_1_0[7] ^ (* src = "crypto_accelerator.v:4050" *) matrix_1_0[4];
  assign _T_1160 = matrix_1_0[6] ^ (* src = "crypto_accelerator.v:4051" *) matrix_1_0[4];
  assign _T_1163 = matrix_1_0[7] ^ (* src = "crypto_accelerator.v:4053" *) matrix_1_0[6];
  assign _T_1166 = matrix_1_0[4] ^ (* src = "crypto_accelerator.v:4055" *) matrix_1_0[3];
  assign _T_1168 = matrix_1_0[3] ^ (* src = "crypto_accelerator.v:4056" *) matrix_1_0[0];
  assign _T_1171 = matrix_1_0[1] ^ (* src = "crypto_accelerator.v:4058" *) matrix_1_0[0];
  assign _T_1173 = matrix_1_0[6] ^ (* src = "crypto_accelerator.v:4059" *) _T_1158;
  assign _T_1176 = _T_1161 ^ (* src = "crypto_accelerator.v:4061" *) _T_1171;
  assign _T_1178 = matrix_1_0[0] ^ (* src = "crypto_accelerator.v:4062" *) _T_1166;
  assign _T_1181 = _T_1164 ^ (* src = "crypto_accelerator.v:4064" *) _T_1169;
  assign _T_1183 = _T_1164 ^ (* src = "crypto_accelerator.v:4065" *) _T_1171;
  assign _T_1185 = _T_1166 ^ (* src = "crypto_accelerator.v:4066" *) _T_1171;
  assign _T_1187 = matrix_1_0[5] ^ (* src = "crypto_accelerator.v:4067" *) _T_1166;
  assign _T_1190 = matrix_1_0[6] ^ (* src = "crypto_accelerator.v:4069" *) matrix_1_0[1];
  assign _T_1192 = matrix_1_0[5] ^ (* src = "crypto_accelerator.v:4070" *) _T_1176;
  assign _T_1195 = _T_1169 ^ (* src = "crypto_accelerator.v:4072" *) _T_1190;
  assign _T_1197 = matrix_1_0[3] ^ (* src = "crypto_accelerator.v:4073" *) _T_1174;
  assign _T_1199 = matrix_1_0[5] ^ (* src = "crypto_accelerator.v:4074" *) matrix_1_0[2];
  assign _T_1202 = matrix_1_0[2] ^ (* src = "crypto_accelerator.v:4076" *) matrix_1_0[1];
  assign _T_1205 = matrix_1_0[5] ^ (* src = "crypto_accelerator.v:4078" *) matrix_1_0[3];
  assign _T_1208 = matrix_1_0[7] ^ (* src = "crypto_accelerator.v:4080" *) _T_1200;
  assign _T_1210 = _T_1161 ^ (* src = "crypto_accelerator.v:4081" *) _T_1200;
  assign _T_1212 = _T_1190 ^ (* src = "crypto_accelerator.v:4082" *) _T_1206;
  assign _T_1214 = _T_1166 ^ (* src = "crypto_accelerator.v:4083" *) _T_1203;
  assign _T_1216 = _T_1181 ^ (* src = "crypto_accelerator.v:4084" *) _T_1214;
  assign _T_1218 = _T_1181 ^ (* src = "crypto_accelerator.v:4085" *) _T_1203;
  assign _T_1220 = _T_1185 ^ (* src = "crypto_accelerator.v:4086" *) _T_1212;
  assign _T_1226 = _T_1218 ^ (* src = "crypto_accelerator.v:4089" *) _T_1222;
  assign _T_1230 = _T_1228 ^ (* src = "crypto_accelerator.v:4091" *) _T_1222;
  assign _T_1236 = _T_1220 ^ (* src = "crypto_accelerator.v:4094" *) _T_1232;
  assign _T_1240 = _T_1238 ^ (* src = "crypto_accelerator.v:4096" *) _T_1232;
  assign _T_1246 = _T_1244 ^ (* src = "crypto_accelerator.v:4099" *) _T_1242;
  assign _T_1250 = _T_1248 ^ (* src = "crypto_accelerator.v:4101" *) _T_1242;
  assign _T_1252 = _T_1226 ^ (* src = "crypto_accelerator.v:4102" *) _T_1224;
  assign _T_1254 = _T_1230 ^ (* src = "crypto_accelerator.v:4103" *) _T_1169;
  assign _T_1256 = _T_1236 ^ (* src = "crypto_accelerator.v:4104" *) _T_1234;
  assign _T_1258 = _T_1240 ^ (* src = "crypto_accelerator.v:4105" *) _T_1250;
  assign _T_1260 = _T_1252 ^ (* src = "crypto_accelerator.v:4106" *) _T_1246;
  assign _T_1262 = _T_1254 ^ (* src = "crypto_accelerator.v:4107" *) _T_1250;
  assign _T_1264 = _T_1256 ^ (* src = "crypto_accelerator.v:4108" *) _T_1246;
  assign _T_1266 = _T_1258 ^ (* src = "crypto_accelerator.v:4109" *) _T_1188;
  assign _T_1268 = _T_1264 ^ (* src = "crypto_accelerator.v:4110" *) _T_1266;
  assign _T_1272 = _T_1262 ^ (* src = "crypto_accelerator.v:4112" *) _T_1270;
  assign _T_1274 = _T_1260 ^ (* src = "crypto_accelerator.v:4113" *) _T_1262;
  assign _T_1276 = _T_1266 ^ (* src = "crypto_accelerator.v:4114" *) _T_1270;
  assign _T_1286 = _T_1274 ^ (* src = "crypto_accelerator.v:4119" *) _T_1270;
  assign _T_1292 = _T_1268 ^ (* src = "crypto_accelerator.v:4122" *) _T_1270;
  assign _T_1294 = _T_1262 ^ (* src = "crypto_accelerator.v:4123" *) _T_1278;
  assign _T_1296 = _T_1284 ^ (* src = "crypto_accelerator.v:4124" *) _T_1286;
  assign _T_1298 = _T_1266 ^ (* src = "crypto_accelerator.v:4125" *) _T_1280;
  assign _T_1300 = _T_1290 ^ (* src = "crypto_accelerator.v:4126" *) _T_1292;
  assign _T_1302 = _T_1296 ^ (* src = "crypto_accelerator.v:4127" *) _T_1300;
  assign _T_1304 = _T_1294 ^ (* src = "crypto_accelerator.v:4128" *) _T_1298;
  assign _T_1306 = _T_1294 ^ (* src = "crypto_accelerator.v:4129" *) _T_1296;
  assign _T_1308 = _T_1298 ^ (* src = "crypto_accelerator.v:4130" *) _T_1300;
  assign _T_1310 = _T_1304 ^ (* src = "crypto_accelerator.v:4131" *) _T_1302;
  assign _T_1348 = _T_1324 ^ (* src = "crypto_accelerator.v:4150" *) _T_1342;
  assign _T_1350 = _T_1336 ^ (* src = "crypto_accelerator.v:4151" *) _T_1338;
  assign _T_1352 = _T_1328 ^ (* src = "crypto_accelerator.v:4152" *) _T_1344;
  assign _T_1354 = _T_1314 ^ (* src = "crypto_accelerator.v:4153" *) _T_1320;
  assign _T_1356 = _T_1316 ^ (* src = "crypto_accelerator.v:4154" *) _T_1332;
  assign _T_1358 = _T_1312 ^ (* src = "crypto_accelerator.v:4155" *) _T_1322;
  assign _T_1360 = _T_1318 ^ (* src = "crypto_accelerator.v:4156" *) _T_1340;
  assign _T_1362 = _T_1348 ^ (* src = "crypto_accelerator.v:4157" *) _T_1350;
  assign _T_1364 = _T_1320 ^ (* src = "crypto_accelerator.v:4158" *) _T_1326;
  assign _T_1366 = _T_1330 ^ (* src = "crypto_accelerator.v:4159" *) _T_1346;
  assign _T_1368 = _T_1334 ^ (* src = "crypto_accelerator.v:4160" *) _T_1356;
  assign _T_1370 = _T_1348 ^ (* src = "crypto_accelerator.v:4161" *) _T_1354;
  assign _T_1372 = _T_1312 ^ (* src = "crypto_accelerator.v:4162" *) _T_1316;
  assign _T_1374 = _T_1318 ^ (* src = "crypto_accelerator.v:4163" *) _T_1322;
  assign _T_1376 = _T_1318 ^ (* src = "crypto_accelerator.v:4164" *) _T_1344;
  assign _T_1378 = _T_1328 ^ (* src = "crypto_accelerator.v:4165" *) _T_1338;
  assign _T_1380 = _T_1334 ^ (* src = "crypto_accelerator.v:4166" *) _T_1342;
  assign _T_1382 = _T_1336 ^ (* src = "crypto_accelerator.v:4167" *) _T_1352;
  assign _T_1384 = _T_1346 ^ (* src = "crypto_accelerator.v:4168" *) _T_1358;
  assign _T_1386 = _T_1352 ^ (* src = "crypto_accelerator.v:4169" *) _T_1354;
  assign _T_1388 = _T_1356 ^ (* src = "crypto_accelerator.v:4170" *) _T_1360;
  assign _T_1390 = _T_1352 ^ (* src = "crypto_accelerator.v:4171" *) _T_1362;
  assign _T_1392 = _T_1362 ^ (* src = "crypto_accelerator.v:4172" *) _T_1364;
  assign _T_1394 = _T_1358 ^ (* src = "crypto_accelerator.v:4173" *) _T_1362;
  assign _T_1396 = _T_1360 ^ (* src = "crypto_accelerator.v:4174" *) _T_1368;
  assign _T_1398 = _T_1366 ^ (* src = "crypto_accelerator.v:4175" *) _T_1370;
  assign _T_1400 = _T_1368 ^ (* src = "crypto_accelerator.v:4176" *) _T_1384;
  assign _T_1402 = _T_1370 ^ (* src = "crypto_accelerator.v:4177" *) _T_1396;
  assign _T_1404 = _T_1378 ^ (* src = "crypto_accelerator.v:4178" *) _T_1388;
  assign _T_1405 = _T_1374 ^ (* src = "crypto_accelerator.v:4179" *) _T_1390;
  assign _T_1406 = _T_1398 ^ (* src = "crypto_accelerator.v:4180" *) _T_1404;
  assign _T_1407 = _T_1382 ^ (* src = "crypto_accelerator.v:4181" *) _T_1402;
  assign _T_1408 = _T_1372 ^ (* src = "crypto_accelerator.v:4182" *) _T_1390;
  assign _T_1409 = _T_1392 ^ (* src = "crypto_accelerator.v:4183" *) _T_1400;
  assign _T_1410 = _T_1386 ^ (* src = "crypto_accelerator.v:4184" *) _T_1394;
  assign _T_1411 = _T_1376 ^ (* src = "crypto_accelerator.v:4185" *) _T_1392;
  assign _T_1412 = _T_1366 ^ (* src = "crypto_accelerator.v:4186" *) _T_1380;
  assign _T_1437 = matrix_0_1[7] ^ (* src = "crypto_accelerator.v:4188" *) matrix_0_1[4];
  assign _T_1439 = matrix_0_1[6] ^ (* src = "crypto_accelerator.v:4189" *) matrix_0_1[4];
  assign _T_1442 = matrix_0_1[7] ^ (* src = "crypto_accelerator.v:4191" *) matrix_0_1[6];
  assign _T_1445 = matrix_0_1[4] ^ (* src = "crypto_accelerator.v:4193" *) matrix_0_1[3];
  assign _T_1447 = matrix_0_1[3] ^ (* src = "crypto_accelerator.v:4194" *) matrix_0_1[0];
  assign _T_1450 = matrix_0_1[1] ^ (* src = "crypto_accelerator.v:4196" *) matrix_0_1[0];
  assign _T_1452 = matrix_0_1[6] ^ (* src = "crypto_accelerator.v:4197" *) _T_1437;
  assign _T_1455 = _T_1440 ^ (* src = "crypto_accelerator.v:4199" *) _T_1450;
  assign _T_1457 = matrix_0_1[0] ^ (* src = "crypto_accelerator.v:4200" *) _T_1445;
  assign _T_1460 = _T_1443 ^ (* src = "crypto_accelerator.v:4202" *) _T_1448;
  assign _T_1462 = _T_1443 ^ (* src = "crypto_accelerator.v:4203" *) _T_1450;
  assign _T_1464 = _T_1445 ^ (* src = "crypto_accelerator.v:4204" *) _T_1450;
  assign _T_1466 = matrix_0_1[5] ^ (* src = "crypto_accelerator.v:4205" *) _T_1445;
  assign _T_1469 = matrix_0_1[6] ^ (* src = "crypto_accelerator.v:4207" *) matrix_0_1[1];
  assign _T_1471 = matrix_0_1[5] ^ (* src = "crypto_accelerator.v:4208" *) _T_1455;
  assign _T_1474 = _T_1448 ^ (* src = "crypto_accelerator.v:4210" *) _T_1469;
  assign _T_1476 = matrix_0_1[3] ^ (* src = "crypto_accelerator.v:4211" *) _T_1453;
  assign _T_1478 = matrix_0_1[5] ^ (* src = "crypto_accelerator.v:4212" *) matrix_0_1[2];
  assign _T_1481 = matrix_0_1[2] ^ (* src = "crypto_accelerator.v:4214" *) matrix_0_1[1];
  assign _T_1484 = matrix_0_1[5] ^ (* src = "crypto_accelerator.v:4216" *) matrix_0_1[3];
  assign _T_1487 = matrix_0_1[7] ^ (* src = "crypto_accelerator.v:4218" *) _T_1479;
  assign _T_1489 = _T_1440 ^ (* src = "crypto_accelerator.v:4219" *) _T_1479;
  assign _T_1491 = _T_1469 ^ (* src = "crypto_accelerator.v:4220" *) _T_1485;
  assign _T_1493 = _T_1445 ^ (* src = "crypto_accelerator.v:4221" *) _T_1482;
  assign _T_1495 = _T_1460 ^ (* src = "crypto_accelerator.v:4222" *) _T_1493;
  assign _T_1497 = _T_1460 ^ (* src = "crypto_accelerator.v:4223" *) _T_1482;
  assign _T_1499 = _T_1464 ^ (* src = "crypto_accelerator.v:4224" *) _T_1491;
  assign _T_1505 = _T_1497 ^ (* src = "crypto_accelerator.v:4227" *) _T_1501;
  assign _T_1509 = _T_1507 ^ (* src = "crypto_accelerator.v:4229" *) _T_1501;
  assign _T_1515 = _T_1499 ^ (* src = "crypto_accelerator.v:4232" *) _T_1511;
  assign _T_1519 = _T_1517 ^ (* src = "crypto_accelerator.v:4234" *) _T_1511;
  assign _T_1525 = _T_1523 ^ (* src = "crypto_accelerator.v:4237" *) _T_1521;
  assign _T_1529 = _T_1527 ^ (* src = "crypto_accelerator.v:4239" *) _T_1521;
  assign _T_1531 = _T_1505 ^ (* src = "crypto_accelerator.v:4240" *) _T_1503;
  assign _T_1533 = _T_1509 ^ (* src = "crypto_accelerator.v:4241" *) _T_1448;
  assign _T_1535 = _T_1515 ^ (* src = "crypto_accelerator.v:4242" *) _T_1513;
  assign _T_1537 = _T_1519 ^ (* src = "crypto_accelerator.v:4243" *) _T_1529;
  assign _T_1539 = _T_1531 ^ (* src = "crypto_accelerator.v:4244" *) _T_1525;
  assign _T_1541 = _T_1533 ^ (* src = "crypto_accelerator.v:4245" *) _T_1529;
  assign _T_1543 = _T_1535 ^ (* src = "crypto_accelerator.v:4246" *) _T_1525;
  assign _T_1545 = _T_1537 ^ (* src = "crypto_accelerator.v:4247" *) _T_1467;
  assign _T_1547 = _T_1543 ^ (* src = "crypto_accelerator.v:4248" *) _T_1545;
  assign _T_1551 = _T_1541 ^ (* src = "crypto_accelerator.v:4250" *) _T_1549;
  assign _T_1553 = _T_1539 ^ (* src = "crypto_accelerator.v:4251" *) _T_1541;
  assign _T_1555 = _T_1545 ^ (* src = "crypto_accelerator.v:4252" *) _T_1549;
  assign _T_1565 = _T_1553 ^ (* src = "crypto_accelerator.v:4257" *) _T_1549;
  assign _T_1571 = _T_1547 ^ (* src = "crypto_accelerator.v:4260" *) _T_1549;
  assign _T_1573 = _T_1541 ^ (* src = "crypto_accelerator.v:4261" *) _T_1557;
  assign _T_1575 = _T_1563 ^ (* src = "crypto_accelerator.v:4262" *) _T_1565;
  assign _T_1577 = _T_1545 ^ (* src = "crypto_accelerator.v:4263" *) _T_1559;
  assign _T_1579 = _T_1569 ^ (* src = "crypto_accelerator.v:4264" *) _T_1571;
  assign _T_1581 = _T_1575 ^ (* src = "crypto_accelerator.v:4265" *) _T_1579;
  assign _T_1583 = _T_1573 ^ (* src = "crypto_accelerator.v:4266" *) _T_1577;
  assign _T_1585 = _T_1573 ^ (* src = "crypto_accelerator.v:4267" *) _T_1575;
  assign _T_1587 = _T_1577 ^ (* src = "crypto_accelerator.v:4268" *) _T_1579;
  assign _T_1589 = _T_1583 ^ (* src = "crypto_accelerator.v:4269" *) _T_1581;
  assign _T_1627 = _T_1603 ^ (* src = "crypto_accelerator.v:4288" *) _T_1621;
  assign _T_1629 = _T_1615 ^ (* src = "crypto_accelerator.v:4289" *) _T_1617;
  assign _T_1631 = _T_1607 ^ (* src = "crypto_accelerator.v:4290" *) _T_1623;
  assign _T_1633 = _T_1593 ^ (* src = "crypto_accelerator.v:4291" *) _T_1599;
  assign _T_1635 = _T_1595 ^ (* src = "crypto_accelerator.v:4292" *) _T_1611;
  assign _T_1637 = _T_1591 ^ (* src = "crypto_accelerator.v:4293" *) _T_1601;
  assign _T_1639 = _T_1597 ^ (* src = "crypto_accelerator.v:4294" *) _T_1619;
  assign _T_1641 = _T_1627 ^ (* src = "crypto_accelerator.v:4295" *) _T_1629;
  assign _T_1643 = _T_1599 ^ (* src = "crypto_accelerator.v:4296" *) _T_1605;
  assign _T_1645 = _T_1609 ^ (* src = "crypto_accelerator.v:4297" *) _T_1625;
  assign _T_1647 = _T_1613 ^ (* src = "crypto_accelerator.v:4298" *) _T_1635;
  assign _T_1649 = _T_1627 ^ (* src = "crypto_accelerator.v:4299" *) _T_1633;
  assign _T_1651 = _T_1591 ^ (* src = "crypto_accelerator.v:4300" *) _T_1595;
  assign _T_1653 = _T_1597 ^ (* src = "crypto_accelerator.v:4301" *) _T_1601;
  assign _T_1655 = _T_1597 ^ (* src = "crypto_accelerator.v:4302" *) _T_1623;
  assign _T_1657 = _T_1607 ^ (* src = "crypto_accelerator.v:4303" *) _T_1617;
  assign _T_1659 = _T_1613 ^ (* src = "crypto_accelerator.v:4304" *) _T_1621;
  assign _T_1661 = _T_1615 ^ (* src = "crypto_accelerator.v:4305" *) _T_1631;
  assign _T_1663 = _T_1625 ^ (* src = "crypto_accelerator.v:4306" *) _T_1637;
  assign _T_1665 = _T_1631 ^ (* src = "crypto_accelerator.v:4307" *) _T_1633;
  assign _T_1667 = _T_1635 ^ (* src = "crypto_accelerator.v:4308" *) _T_1639;
  assign _T_1669 = _T_1631 ^ (* src = "crypto_accelerator.v:4309" *) _T_1641;
  assign _T_1671 = _T_1641 ^ (* src = "crypto_accelerator.v:4310" *) _T_1643;
  assign _T_1673 = _T_1637 ^ (* src = "crypto_accelerator.v:4311" *) _T_1641;
  assign _T_1675 = _T_1639 ^ (* src = "crypto_accelerator.v:4312" *) _T_1647;
  assign _T_1677 = _T_1645 ^ (* src = "crypto_accelerator.v:4313" *) _T_1649;
  assign _T_1679 = _T_1647 ^ (* src = "crypto_accelerator.v:4314" *) _T_1663;
  assign _T_1681 = _T_1649 ^ (* src = "crypto_accelerator.v:4315" *) _T_1675;
  assign _T_1683 = _T_1657 ^ (* src = "crypto_accelerator.v:4316" *) _T_1667;
  assign _T_1684 = _T_1653 ^ (* src = "crypto_accelerator.v:4317" *) _T_1669;
  assign _T_1685 = _T_1677 ^ (* src = "crypto_accelerator.v:4318" *) _T_1683;
  assign _T_1686 = _T_1661 ^ (* src = "crypto_accelerator.v:4319" *) _T_1681;
  assign _T_1687 = _T_1651 ^ (* src = "crypto_accelerator.v:4320" *) _T_1669;
  assign _T_1688 = _T_1671 ^ (* src = "crypto_accelerator.v:4321" *) _T_1679;
  assign _T_1689 = _T_1665 ^ (* src = "crypto_accelerator.v:4322" *) _T_1673;
  assign _T_1690 = _T_1655 ^ (* src = "crypto_accelerator.v:4323" *) _T_1671;
  assign _T_1691 = _T_1645 ^ (* src = "crypto_accelerator.v:4324" *) _T_1659;
  assign _T_1716 = matrix_3_2[7] ^ (* src = "crypto_accelerator.v:4326" *) matrix_3_2[4];
  assign _T_1718 = matrix_3_2[6] ^ (* src = "crypto_accelerator.v:4327" *) matrix_3_2[4];
  assign _T_1721 = matrix_3_2[7] ^ (* src = "crypto_accelerator.v:4329" *) matrix_3_2[6];
  assign _T_1724 = matrix_3_2[4] ^ (* src = "crypto_accelerator.v:4331" *) matrix_3_2[3];
  assign _T_1726 = matrix_3_2[3] ^ (* src = "crypto_accelerator.v:4332" *) matrix_3_2[0];
  assign _T_1729 = matrix_3_2[1] ^ (* src = "crypto_accelerator.v:4334" *) matrix_3_2[0];
  assign _T_1731 = matrix_3_2[6] ^ (* src = "crypto_accelerator.v:4335" *) _T_1716;
  assign _T_1734 = _T_1719 ^ (* src = "crypto_accelerator.v:4337" *) _T_1729;
  assign _T_1736 = matrix_3_2[0] ^ (* src = "crypto_accelerator.v:4338" *) _T_1724;
  assign _T_1739 = _T_1722 ^ (* src = "crypto_accelerator.v:4340" *) _T_1727;
  assign _T_1741 = _T_1722 ^ (* src = "crypto_accelerator.v:4341" *) _T_1729;
  assign _T_1743 = _T_1724 ^ (* src = "crypto_accelerator.v:4342" *) _T_1729;
  assign _T_1745 = matrix_3_2[5] ^ (* src = "crypto_accelerator.v:4343" *) _T_1724;
  assign _T_1748 = matrix_3_2[6] ^ (* src = "crypto_accelerator.v:4345" *) matrix_3_2[1];
  assign _T_1750 = matrix_3_2[5] ^ (* src = "crypto_accelerator.v:4346" *) _T_1734;
  assign _T_1753 = _T_1727 ^ (* src = "crypto_accelerator.v:4348" *) _T_1748;
  assign _T_1755 = matrix_3_2[3] ^ (* src = "crypto_accelerator.v:4349" *) _T_1732;
  assign _T_1757 = matrix_3_2[5] ^ (* src = "crypto_accelerator.v:4350" *) matrix_3_2[2];
  assign _T_1760 = matrix_3_2[2] ^ (* src = "crypto_accelerator.v:4352" *) matrix_3_2[1];
  assign _T_1763 = matrix_3_2[5] ^ (* src = "crypto_accelerator.v:4354" *) matrix_3_2[3];
  assign _T_1766 = matrix_3_2[7] ^ (* src = "crypto_accelerator.v:4356" *) _T_1758;
  assign _T_1768 = _T_1719 ^ (* src = "crypto_accelerator.v:4357" *) _T_1758;
  assign _T_1770 = _T_1748 ^ (* src = "crypto_accelerator.v:4358" *) _T_1764;
  assign _T_1772 = _T_1724 ^ (* src = "crypto_accelerator.v:4359" *) _T_1761;
  assign _T_1774 = _T_1739 ^ (* src = "crypto_accelerator.v:4360" *) _T_1772;
  assign _T_1776 = _T_1739 ^ (* src = "crypto_accelerator.v:4361" *) _T_1761;
  assign _T_1778 = _T_1743 ^ (* src = "crypto_accelerator.v:4362" *) _T_1770;
  assign _T_1784 = _T_1776 ^ (* src = "crypto_accelerator.v:4365" *) _T_1780;
  assign _T_1788 = _T_1786 ^ (* src = "crypto_accelerator.v:4367" *) _T_1780;
  assign _T_1794 = _T_1778 ^ (* src = "crypto_accelerator.v:4370" *) _T_1790;
  assign _T_1798 = _T_1796 ^ (* src = "crypto_accelerator.v:4372" *) _T_1790;
  assign _T_1804 = _T_1802 ^ (* src = "crypto_accelerator.v:4375" *) _T_1800;
  assign _T_1808 = _T_1806 ^ (* src = "crypto_accelerator.v:4377" *) _T_1800;
  assign _T_1810 = _T_1784 ^ (* src = "crypto_accelerator.v:4378" *) _T_1782;
  assign _T_1812 = _T_1788 ^ (* src = "crypto_accelerator.v:4379" *) _T_1727;
  assign _T_1814 = _T_1794 ^ (* src = "crypto_accelerator.v:4380" *) _T_1792;
  assign _T_1816 = _T_1798 ^ (* src = "crypto_accelerator.v:4381" *) _T_1808;
  assign _T_1818 = _T_1810 ^ (* src = "crypto_accelerator.v:4382" *) _T_1804;
  assign _T_1820 = _T_1812 ^ (* src = "crypto_accelerator.v:4383" *) _T_1808;
  assign _T_1822 = _T_1814 ^ (* src = "crypto_accelerator.v:4384" *) _T_1804;
  assign _T_1824 = _T_1816 ^ (* src = "crypto_accelerator.v:4385" *) _T_1746;
  assign _T_1826 = _T_1822 ^ (* src = "crypto_accelerator.v:4386" *) _T_1824;
  assign _T_1830 = _T_1820 ^ (* src = "crypto_accelerator.v:4388" *) _T_1828;
  assign _T_1832 = _T_1818 ^ (* src = "crypto_accelerator.v:4389" *) _T_1820;
  assign _T_1834 = _T_1824 ^ (* src = "crypto_accelerator.v:4390" *) _T_1828;
  assign _T_1844 = _T_1832 ^ (* src = "crypto_accelerator.v:4395" *) _T_1828;
  assign _T_1850 = _T_1826 ^ (* src = "crypto_accelerator.v:4398" *) _T_1828;
  assign _T_1852 = _T_1820 ^ (* src = "crypto_accelerator.v:4399" *) _T_1836;
  assign _T_1854 = _T_1842 ^ (* src = "crypto_accelerator.v:4400" *) _T_1844;
  assign _T_1856 = _T_1824 ^ (* src = "crypto_accelerator.v:4401" *) _T_1838;
  assign _T_1858 = _T_1848 ^ (* src = "crypto_accelerator.v:4402" *) _T_1850;
  assign _T_1860 = _T_1854 ^ (* src = "crypto_accelerator.v:4403" *) _T_1858;
  assign _T_1862 = _T_1852 ^ (* src = "crypto_accelerator.v:4404" *) _T_1856;
  assign _T_1864 = _T_1852 ^ (* src = "crypto_accelerator.v:4405" *) _T_1854;
  assign _T_1866 = _T_1856 ^ (* src = "crypto_accelerator.v:4406" *) _T_1858;
  assign _T_1868 = _T_1862 ^ (* src = "crypto_accelerator.v:4407" *) _T_1860;
  assign _T_1906 = _T_1882 ^ (* src = "crypto_accelerator.v:4426" *) _T_1900;
  assign _T_1908 = _T_1894 ^ (* src = "crypto_accelerator.v:4427" *) _T_1896;
  assign _T_1910 = _T_1886 ^ (* src = "crypto_accelerator.v:4428" *) _T_1902;
  assign _T_1912 = _T_1872 ^ (* src = "crypto_accelerator.v:4429" *) _T_1878;
  assign _T_1914 = _T_1874 ^ (* src = "crypto_accelerator.v:4430" *) _T_1890;
  assign _T_1916 = _T_1870 ^ (* src = "crypto_accelerator.v:4431" *) _T_1880;
  assign _T_1918 = _T_1876 ^ (* src = "crypto_accelerator.v:4432" *) _T_1898;
  assign _T_1920 = _T_1906 ^ (* src = "crypto_accelerator.v:4433" *) _T_1908;
  assign _T_1922 = _T_1878 ^ (* src = "crypto_accelerator.v:4434" *) _T_1884;
  assign _T_1924 = _T_1888 ^ (* src = "crypto_accelerator.v:4435" *) _T_1904;
  assign _T_1926 = _T_1892 ^ (* src = "crypto_accelerator.v:4436" *) _T_1914;
  assign _T_1928 = _T_1906 ^ (* src = "crypto_accelerator.v:4437" *) _T_1912;
  assign _T_1930 = _T_1870 ^ (* src = "crypto_accelerator.v:4438" *) _T_1874;
  assign _T_1932 = _T_1876 ^ (* src = "crypto_accelerator.v:4439" *) _T_1880;
  assign _T_1934 = _T_1876 ^ (* src = "crypto_accelerator.v:4440" *) _T_1902;
  assign _T_1936 = _T_1886 ^ (* src = "crypto_accelerator.v:4441" *) _T_1896;
  assign _T_1938 = _T_1892 ^ (* src = "crypto_accelerator.v:4442" *) _T_1900;
  assign _T_1940 = _T_1894 ^ (* src = "crypto_accelerator.v:4443" *) _T_1910;
  assign _T_1942 = _T_1904 ^ (* src = "crypto_accelerator.v:4444" *) _T_1916;
  assign _T_1944 = _T_1910 ^ (* src = "crypto_accelerator.v:4445" *) _T_1912;
  assign _T_1946 = _T_1914 ^ (* src = "crypto_accelerator.v:4446" *) _T_1918;
  assign _T_1948 = _T_1910 ^ (* src = "crypto_accelerator.v:4447" *) _T_1920;
  assign _T_1950 = _T_1920 ^ (* src = "crypto_accelerator.v:4448" *) _T_1922;
  assign _T_1952 = _T_1916 ^ (* src = "crypto_accelerator.v:4449" *) _T_1920;
  assign _T_1954 = _T_1918 ^ (* src = "crypto_accelerator.v:4450" *) _T_1926;
  assign _T_1956 = _T_1924 ^ (* src = "crypto_accelerator.v:4451" *) _T_1928;
  assign _T_1958 = _T_1926 ^ (* src = "crypto_accelerator.v:4452" *) _T_1942;
  assign _T_1960 = _T_1928 ^ (* src = "crypto_accelerator.v:4453" *) _T_1954;
  assign _T_1962 = _T_1936 ^ (* src = "crypto_accelerator.v:4454" *) _T_1946;
  assign _T_1963 = _T_1932 ^ (* src = "crypto_accelerator.v:4455" *) _T_1948;
  assign _T_1964 = _T_1956 ^ (* src = "crypto_accelerator.v:4456" *) _T_1962;
  assign _T_1965 = _T_1940 ^ (* src = "crypto_accelerator.v:4457" *) _T_1960;
  assign _T_1966 = _T_1930 ^ (* src = "crypto_accelerator.v:4458" *) _T_1948;
  assign _T_1967 = _T_1950 ^ (* src = "crypto_accelerator.v:4459" *) _T_1958;
  assign _T_1968 = _T_1944 ^ (* src = "crypto_accelerator.v:4460" *) _T_1952;
  assign _T_1969 = _T_1934 ^ (* src = "crypto_accelerator.v:4461" *) _T_1950;
  assign _T_1970 = _T_1924 ^ (* src = "crypto_accelerator.v:4462" *) _T_1938;
  assign _T_1995 = matrix_2_3[7] ^ (* src = "crypto_accelerator.v:4464" *) matrix_2_3[4];
  assign _T_1997 = matrix_2_3[6] ^ (* src = "crypto_accelerator.v:4465" *) matrix_2_3[4];
  assign _T_2000 = matrix_2_3[7] ^ (* src = "crypto_accelerator.v:4467" *) matrix_2_3[6];
  assign _T_2003 = matrix_2_3[4] ^ (* src = "crypto_accelerator.v:4469" *) matrix_2_3[3];
  assign _T_2005 = matrix_2_3[3] ^ (* src = "crypto_accelerator.v:4470" *) matrix_2_3[0];
  assign _T_2008 = matrix_2_3[1] ^ (* src = "crypto_accelerator.v:4472" *) matrix_2_3[0];
  assign _T_2010 = matrix_2_3[6] ^ (* src = "crypto_accelerator.v:4473" *) _T_1995;
  assign _T_2013 = _T_1998 ^ (* src = "crypto_accelerator.v:4475" *) _T_2008;
  assign _T_2015 = matrix_2_3[0] ^ (* src = "crypto_accelerator.v:4476" *) _T_2003;
  assign _T_2018 = _T_2001 ^ (* src = "crypto_accelerator.v:4478" *) _T_2006;
  assign _T_2020 = _T_2001 ^ (* src = "crypto_accelerator.v:4479" *) _T_2008;
  assign _T_2022 = _T_2003 ^ (* src = "crypto_accelerator.v:4480" *) _T_2008;
  assign _T_2024 = matrix_2_3[5] ^ (* src = "crypto_accelerator.v:4481" *) _T_2003;
  assign _T_2027 = matrix_2_3[6] ^ (* src = "crypto_accelerator.v:4483" *) matrix_2_3[1];
  assign _T_2029 = matrix_2_3[5] ^ (* src = "crypto_accelerator.v:4484" *) _T_2013;
  assign _T_2032 = _T_2006 ^ (* src = "crypto_accelerator.v:4486" *) _T_2027;
  assign _T_2034 = matrix_2_3[3] ^ (* src = "crypto_accelerator.v:4487" *) _T_2011;
  assign _T_2036 = matrix_2_3[5] ^ (* src = "crypto_accelerator.v:4488" *) matrix_2_3[2];
  assign _T_2039 = matrix_2_3[2] ^ (* src = "crypto_accelerator.v:4490" *) matrix_2_3[1];
  assign _T_2042 = matrix_2_3[5] ^ (* src = "crypto_accelerator.v:4492" *) matrix_2_3[3];
  assign _T_2045 = matrix_2_3[7] ^ (* src = "crypto_accelerator.v:4494" *) _T_2037;
  assign _T_2047 = _T_1998 ^ (* src = "crypto_accelerator.v:4495" *) _T_2037;
  assign _T_2049 = _T_2027 ^ (* src = "crypto_accelerator.v:4496" *) _T_2043;
  assign _T_2051 = _T_2003 ^ (* src = "crypto_accelerator.v:4497" *) _T_2040;
  assign _T_2053 = _T_2018 ^ (* src = "crypto_accelerator.v:4498" *) _T_2051;
  assign _T_2055 = _T_2018 ^ (* src = "crypto_accelerator.v:4499" *) _T_2040;
  assign _T_2057 = _T_2022 ^ (* src = "crypto_accelerator.v:4500" *) _T_2049;
  assign _T_2063 = _T_2055 ^ (* src = "crypto_accelerator.v:4503" *) _T_2059;
  assign _T_2067 = _T_2065 ^ (* src = "crypto_accelerator.v:4505" *) _T_2059;
  assign _T_2073 = _T_2057 ^ (* src = "crypto_accelerator.v:4508" *) _T_2069;
  assign _T_2077 = _T_2075 ^ (* src = "crypto_accelerator.v:4510" *) _T_2069;
  assign _T_2083 = _T_2081 ^ (* src = "crypto_accelerator.v:4513" *) _T_2079;
  assign _T_2087 = _T_2085 ^ (* src = "crypto_accelerator.v:4515" *) _T_2079;
  assign _T_2089 = _T_2063 ^ (* src = "crypto_accelerator.v:4516" *) _T_2061;
  assign _T_2091 = _T_2067 ^ (* src = "crypto_accelerator.v:4517" *) _T_2006;
  assign _T_2093 = _T_2073 ^ (* src = "crypto_accelerator.v:4518" *) _T_2071;
  assign _T_2095 = _T_2077 ^ (* src = "crypto_accelerator.v:4519" *) _T_2087;
  assign _T_2097 = _T_2089 ^ (* src = "crypto_accelerator.v:4520" *) _T_2083;
  assign _T_2099 = _T_2091 ^ (* src = "crypto_accelerator.v:4521" *) _T_2087;
  assign _T_2101 = _T_2093 ^ (* src = "crypto_accelerator.v:4522" *) _T_2083;
  assign _T_2103 = _T_2095 ^ (* src = "crypto_accelerator.v:4523" *) _T_2025;
  assign _T_2105 = _T_2101 ^ (* src = "crypto_accelerator.v:4524" *) _T_2103;
  assign _T_2109 = _T_2099 ^ (* src = "crypto_accelerator.v:4526" *) _T_2107;
  assign _T_2111 = _T_2097 ^ (* src = "crypto_accelerator.v:4527" *) _T_2099;
  assign _T_2113 = _T_2103 ^ (* src = "crypto_accelerator.v:4528" *) _T_2107;
  assign _T_2123 = _T_2111 ^ (* src = "crypto_accelerator.v:4533" *) _T_2107;
  assign _T_2129 = _T_2105 ^ (* src = "crypto_accelerator.v:4536" *) _T_2107;
  assign _T_2131 = _T_2099 ^ (* src = "crypto_accelerator.v:4537" *) _T_2115;
  assign _T_2133 = _T_2121 ^ (* src = "crypto_accelerator.v:4538" *) _T_2123;
  assign _T_2135 = _T_2103 ^ (* src = "crypto_accelerator.v:4539" *) _T_2117;
  assign _T_2137 = _T_2127 ^ (* src = "crypto_accelerator.v:4540" *) _T_2129;
  assign _T_2139 = _T_2133 ^ (* src = "crypto_accelerator.v:4541" *) _T_2137;
  assign _T_2141 = _T_2131 ^ (* src = "crypto_accelerator.v:4542" *) _T_2135;
  assign _T_2143 = _T_2131 ^ (* src = "crypto_accelerator.v:4543" *) _T_2133;
  assign _T_2145 = _T_2135 ^ (* src = "crypto_accelerator.v:4544" *) _T_2137;
  assign _T_2147 = _T_2141 ^ (* src = "crypto_accelerator.v:4545" *) _T_2139;
  assign _T_2185 = _T_2161 ^ (* src = "crypto_accelerator.v:4564" *) _T_2179;
  assign _T_2187 = _T_2173 ^ (* src = "crypto_accelerator.v:4565" *) _T_2175;
  assign _T_2189 = _T_2165 ^ (* src = "crypto_accelerator.v:4566" *) _T_2181;
  assign _T_2191 = _T_2151 ^ (* src = "crypto_accelerator.v:4567" *) _T_2157;
  assign _T_2193 = _T_2153 ^ (* src = "crypto_accelerator.v:4568" *) _T_2169;
  assign _T_2195 = _T_2149 ^ (* src = "crypto_accelerator.v:4569" *) _T_2159;
  assign _T_2197 = _T_2155 ^ (* src = "crypto_accelerator.v:4570" *) _T_2177;
  assign _T_2199 = _T_2185 ^ (* src = "crypto_accelerator.v:4571" *) _T_2187;
  assign _T_2201 = _T_2157 ^ (* src = "crypto_accelerator.v:4572" *) _T_2163;
  assign _T_2203 = _T_2167 ^ (* src = "crypto_accelerator.v:4573" *) _T_2183;
  assign _T_2205 = _T_2171 ^ (* src = "crypto_accelerator.v:4574" *) _T_2193;
  assign _T_2207 = _T_2185 ^ (* src = "crypto_accelerator.v:4575" *) _T_2191;
  assign _T_2209 = _T_2149 ^ (* src = "crypto_accelerator.v:4576" *) _T_2153;
  assign _T_2211 = _T_2155 ^ (* src = "crypto_accelerator.v:4577" *) _T_2159;
  assign _T_2213 = _T_2155 ^ (* src = "crypto_accelerator.v:4578" *) _T_2181;
  assign _T_2215 = _T_2165 ^ (* src = "crypto_accelerator.v:4579" *) _T_2175;
  assign _T_2217 = _T_2171 ^ (* src = "crypto_accelerator.v:4580" *) _T_2179;
  assign _T_2219 = _T_2173 ^ (* src = "crypto_accelerator.v:4581" *) _T_2189;
  assign _T_2221 = _T_2183 ^ (* src = "crypto_accelerator.v:4582" *) _T_2195;
  assign _T_2223 = _T_2189 ^ (* src = "crypto_accelerator.v:4583" *) _T_2191;
  assign _T_2225 = _T_2193 ^ (* src = "crypto_accelerator.v:4584" *) _T_2197;
  assign _T_2227 = _T_2189 ^ (* src = "crypto_accelerator.v:4585" *) _T_2199;
  assign _T_2229 = _T_2199 ^ (* src = "crypto_accelerator.v:4586" *) _T_2201;
  assign _T_2231 = _T_2195 ^ (* src = "crypto_accelerator.v:4587" *) _T_2199;
  assign _T_2233 = _T_2197 ^ (* src = "crypto_accelerator.v:4588" *) _T_2205;
  assign _T_2235 = _T_2203 ^ (* src = "crypto_accelerator.v:4589" *) _T_2207;
  assign _T_2237 = _T_2205 ^ (* src = "crypto_accelerator.v:4590" *) _T_2221;
  assign _T_2239 = _T_2207 ^ (* src = "crypto_accelerator.v:4591" *) _T_2233;
  assign _T_2241 = _T_2215 ^ (* src = "crypto_accelerator.v:4592" *) _T_2225;
  assign _T_2242 = _T_2211 ^ (* src = "crypto_accelerator.v:4593" *) _T_2227;
  assign _T_2243 = _T_2235 ^ (* src = "crypto_accelerator.v:4594" *) _T_2241;
  assign _T_2244 = _T_2219 ^ (* src = "crypto_accelerator.v:4595" *) _T_2239;
  assign _T_2245 = _T_2209 ^ (* src = "crypto_accelerator.v:4596" *) _T_2227;
  assign _T_2246 = _T_2229 ^ (* src = "crypto_accelerator.v:4597" *) _T_2237;
  assign _T_2247 = _T_2223 ^ (* src = "crypto_accelerator.v:4598" *) _T_2231;
  assign _T_2248 = _T_2213 ^ (* src = "crypto_accelerator.v:4599" *) _T_2229;
  assign _T_2249 = _T_2203 ^ (* src = "crypto_accelerator.v:4600" *) _T_2217;
  assign _T_2275 = matrix_2_0[7] ^ (* src = "crypto_accelerator.v:4602" *) matrix_2_0[4];
  assign _T_2277 = matrix_2_0[6] ^ (* src = "crypto_accelerator.v:4603" *) matrix_2_0[4];
  assign _T_2280 = matrix_2_0[7] ^ (* src = "crypto_accelerator.v:4605" *) matrix_2_0[6];
  assign _T_2283 = matrix_2_0[4] ^ (* src = "crypto_accelerator.v:4607" *) matrix_2_0[3];
  assign _T_2285 = matrix_2_0[3] ^ (* src = "crypto_accelerator.v:4608" *) matrix_2_0[0];
  assign _T_2288 = matrix_2_0[1] ^ (* src = "crypto_accelerator.v:4610" *) matrix_2_0[0];
  assign _T_2290 = matrix_2_0[6] ^ (* src = "crypto_accelerator.v:4611" *) _T_2275;
  assign _T_2293 = _T_2278 ^ (* src = "crypto_accelerator.v:4613" *) _T_2288;
  assign _T_2295 = matrix_2_0[0] ^ (* src = "crypto_accelerator.v:4614" *) _T_2283;
  assign _T_2298 = _T_2281 ^ (* src = "crypto_accelerator.v:4616" *) _T_2286;
  assign _T_2300 = _T_2281 ^ (* src = "crypto_accelerator.v:4617" *) _T_2288;
  assign _T_2302 = _T_2283 ^ (* src = "crypto_accelerator.v:4618" *) _T_2288;
  assign _T_2304 = matrix_2_0[5] ^ (* src = "crypto_accelerator.v:4619" *) _T_2283;
  assign _T_2307 = matrix_2_0[6] ^ (* src = "crypto_accelerator.v:4621" *) matrix_2_0[1];
  assign _T_2309 = matrix_2_0[5] ^ (* src = "crypto_accelerator.v:4622" *) _T_2293;
  assign _T_2312 = _T_2286 ^ (* src = "crypto_accelerator.v:4624" *) _T_2307;
  assign _T_2314 = matrix_2_0[3] ^ (* src = "crypto_accelerator.v:4625" *) _T_2291;
  assign _T_2316 = matrix_2_0[5] ^ (* src = "crypto_accelerator.v:4626" *) matrix_2_0[2];
  assign _T_2319 = matrix_2_0[2] ^ (* src = "crypto_accelerator.v:4628" *) matrix_2_0[1];
  assign _T_2322 = matrix_2_0[5] ^ (* src = "crypto_accelerator.v:4630" *) matrix_2_0[3];
  assign _T_2325 = matrix_2_0[7] ^ (* src = "crypto_accelerator.v:4632" *) _T_2317;
  assign _T_2327 = _T_2278 ^ (* src = "crypto_accelerator.v:4633" *) _T_2317;
  assign _T_2329 = _T_2307 ^ (* src = "crypto_accelerator.v:4634" *) _T_2323;
  assign _T_2331 = _T_2283 ^ (* src = "crypto_accelerator.v:4635" *) _T_2320;
  assign _T_2333 = _T_2298 ^ (* src = "crypto_accelerator.v:4636" *) _T_2331;
  assign _T_2335 = _T_2298 ^ (* src = "crypto_accelerator.v:4637" *) _T_2320;
  assign _T_2337 = _T_2302 ^ (* src = "crypto_accelerator.v:4638" *) _T_2329;
  assign _T_2343 = _T_2335 ^ (* src = "crypto_accelerator.v:4641" *) _T_2339;
  assign _T_2347 = _T_2345 ^ (* src = "crypto_accelerator.v:4643" *) _T_2339;
  assign _T_2353 = _T_2337 ^ (* src = "crypto_accelerator.v:4646" *) _T_2349;
  assign _T_2357 = _T_2355 ^ (* src = "crypto_accelerator.v:4648" *) _T_2349;
  assign _T_2363 = _T_2361 ^ (* src = "crypto_accelerator.v:4651" *) _T_2359;
  assign _T_2367 = _T_2365 ^ (* src = "crypto_accelerator.v:4653" *) _T_2359;
  assign _T_2369 = _T_2343 ^ (* src = "crypto_accelerator.v:4654" *) _T_2341;
  assign _T_2371 = _T_2347 ^ (* src = "crypto_accelerator.v:4655" *) _T_2286;
  assign _T_2373 = _T_2353 ^ (* src = "crypto_accelerator.v:4656" *) _T_2351;
  assign _T_2375 = _T_2357 ^ (* src = "crypto_accelerator.v:4657" *) _T_2367;
  assign _T_2377 = _T_2369 ^ (* src = "crypto_accelerator.v:4658" *) _T_2363;
  assign _T_2379 = _T_2371 ^ (* src = "crypto_accelerator.v:4659" *) _T_2367;
  assign _T_2381 = _T_2373 ^ (* src = "crypto_accelerator.v:4660" *) _T_2363;
  assign _T_2383 = _T_2375 ^ (* src = "crypto_accelerator.v:4661" *) _T_2305;
  assign _T_2385 = _T_2381 ^ (* src = "crypto_accelerator.v:4662" *) _T_2383;
  assign _T_2389 = _T_2379 ^ (* src = "crypto_accelerator.v:4664" *) _T_2387;
  assign _T_2391 = _T_2377 ^ (* src = "crypto_accelerator.v:4665" *) _T_2379;
  assign _T_2393 = _T_2383 ^ (* src = "crypto_accelerator.v:4666" *) _T_2387;
  assign _T_2403 = _T_2391 ^ (* src = "crypto_accelerator.v:4671" *) _T_2387;
  assign _T_2409 = _T_2385 ^ (* src = "crypto_accelerator.v:4674" *) _T_2387;
  assign _T_2411 = _T_2379 ^ (* src = "crypto_accelerator.v:4675" *) _T_2395;
  assign _T_2413 = _T_2401 ^ (* src = "crypto_accelerator.v:4676" *) _T_2403;
  assign _T_2415 = _T_2383 ^ (* src = "crypto_accelerator.v:4677" *) _T_2397;
  assign _T_2417 = _T_2407 ^ (* src = "crypto_accelerator.v:4678" *) _T_2409;
  assign _T_2419 = _T_2413 ^ (* src = "crypto_accelerator.v:4679" *) _T_2417;
  assign _T_2421 = _T_2411 ^ (* src = "crypto_accelerator.v:4680" *) _T_2415;
  assign _T_2423 = _T_2411 ^ (* src = "crypto_accelerator.v:4681" *) _T_2413;
  assign _T_2425 = _T_2415 ^ (* src = "crypto_accelerator.v:4682" *) _T_2417;
  assign _T_2427 = _T_2421 ^ (* src = "crypto_accelerator.v:4683" *) _T_2419;
  assign _T_2465 = _T_2441 ^ (* src = "crypto_accelerator.v:4702" *) _T_2459;
  assign _T_2467 = _T_2453 ^ (* src = "crypto_accelerator.v:4703" *) _T_2455;
  assign _T_2469 = _T_2445 ^ (* src = "crypto_accelerator.v:4704" *) _T_2461;
  assign _T_2471 = _T_2431 ^ (* src = "crypto_accelerator.v:4705" *) _T_2437;
  assign _T_2473 = _T_2433 ^ (* src = "crypto_accelerator.v:4706" *) _T_2449;
  assign _T_2475 = _T_2429 ^ (* src = "crypto_accelerator.v:4707" *) _T_2439;
  assign _T_2477 = _T_2435 ^ (* src = "crypto_accelerator.v:4708" *) _T_2457;
  assign _T_2479 = _T_2465 ^ (* src = "crypto_accelerator.v:4709" *) _T_2467;
  assign _T_2481 = _T_2437 ^ (* src = "crypto_accelerator.v:4710" *) _T_2443;
  assign _T_2483 = _T_2447 ^ (* src = "crypto_accelerator.v:4711" *) _T_2463;
  assign _T_2485 = _T_2451 ^ (* src = "crypto_accelerator.v:4712" *) _T_2473;
  assign _T_2487 = _T_2465 ^ (* src = "crypto_accelerator.v:4713" *) _T_2471;
  assign _T_2489 = _T_2429 ^ (* src = "crypto_accelerator.v:4714" *) _T_2433;
  assign _T_2491 = _T_2435 ^ (* src = "crypto_accelerator.v:4715" *) _T_2439;
  assign _T_2493 = _T_2435 ^ (* src = "crypto_accelerator.v:4716" *) _T_2461;
  assign _T_2495 = _T_2445 ^ (* src = "crypto_accelerator.v:4717" *) _T_2455;
  assign _T_2497 = _T_2451 ^ (* src = "crypto_accelerator.v:4718" *) _T_2459;
  assign _T_2499 = _T_2453 ^ (* src = "crypto_accelerator.v:4719" *) _T_2469;
  assign _T_2501 = _T_2463 ^ (* src = "crypto_accelerator.v:4720" *) _T_2475;
  assign _T_2503 = _T_2469 ^ (* src = "crypto_accelerator.v:4721" *) _T_2471;
  assign _T_2505 = _T_2473 ^ (* src = "crypto_accelerator.v:4722" *) _T_2477;
  assign _T_2507 = _T_2469 ^ (* src = "crypto_accelerator.v:4723" *) _T_2479;
  assign _T_2509 = _T_2479 ^ (* src = "crypto_accelerator.v:4724" *) _T_2481;
  assign _T_2511 = _T_2475 ^ (* src = "crypto_accelerator.v:4725" *) _T_2479;
  assign _T_2513 = _T_2477 ^ (* src = "crypto_accelerator.v:4726" *) _T_2485;
  assign _T_2515 = _T_2483 ^ (* src = "crypto_accelerator.v:4727" *) _T_2487;
  assign _T_2517 = _T_2485 ^ (* src = "crypto_accelerator.v:4728" *) _T_2501;
  assign _T_2519 = _T_2487 ^ (* src = "crypto_accelerator.v:4729" *) _T_2513;
  assign _T_2521 = _T_2495 ^ (* src = "crypto_accelerator.v:4730" *) _T_2505;
  assign _T_2522 = _T_2491 ^ (* src = "crypto_accelerator.v:4731" *) _T_2507;
  assign _T_2523 = _T_2515 ^ (* src = "crypto_accelerator.v:4732" *) _T_2521;
  assign _T_2524 = _T_2499 ^ (* src = "crypto_accelerator.v:4733" *) _T_2519;
  assign _T_2525 = _T_2489 ^ (* src = "crypto_accelerator.v:4734" *) _T_2507;
  assign _T_2526 = _T_2509 ^ (* src = "crypto_accelerator.v:4735" *) _T_2517;
  assign _T_2527 = _T_2503 ^ (* src = "crypto_accelerator.v:4736" *) _T_2511;
  assign _T_2528 = _T_2493 ^ (* src = "crypto_accelerator.v:4737" *) _T_2509;
  assign _T_2529 = _T_2483 ^ (* src = "crypto_accelerator.v:4738" *) _T_2497;
  assign _T_2554 = matrix_1_1[7] ^ (* src = "crypto_accelerator.v:4740" *) matrix_1_1[4];
  assign _T_2556 = matrix_1_1[6] ^ (* src = "crypto_accelerator.v:4741" *) matrix_1_1[4];
  assign _T_2559 = matrix_1_1[7] ^ (* src = "crypto_accelerator.v:4743" *) matrix_1_1[6];
  assign _T_2562 = matrix_1_1[4] ^ (* src = "crypto_accelerator.v:4745" *) matrix_1_1[3];
  assign _T_2564 = matrix_1_1[3] ^ (* src = "crypto_accelerator.v:4746" *) matrix_1_1[0];
  assign _T_2567 = matrix_1_1[1] ^ (* src = "crypto_accelerator.v:4748" *) matrix_1_1[0];
  assign _T_2569 = matrix_1_1[6] ^ (* src = "crypto_accelerator.v:4749" *) _T_2554;
  assign _T_2572 = _T_2557 ^ (* src = "crypto_accelerator.v:4751" *) _T_2567;
  assign _T_2574 = matrix_1_1[0] ^ (* src = "crypto_accelerator.v:4752" *) _T_2562;
  assign _T_2577 = _T_2560 ^ (* src = "crypto_accelerator.v:4754" *) _T_2565;
  assign _T_2579 = _T_2560 ^ (* src = "crypto_accelerator.v:4755" *) _T_2567;
  assign _T_2581 = _T_2562 ^ (* src = "crypto_accelerator.v:4756" *) _T_2567;
  assign _T_2583 = matrix_1_1[5] ^ (* src = "crypto_accelerator.v:4757" *) _T_2562;
  assign _T_2586 = matrix_1_1[6] ^ (* src = "crypto_accelerator.v:4759" *) matrix_1_1[1];
  assign _T_2588 = matrix_1_1[5] ^ (* src = "crypto_accelerator.v:4760" *) _T_2572;
  assign _T_2591 = _T_2565 ^ (* src = "crypto_accelerator.v:4762" *) _T_2586;
  assign _T_2593 = matrix_1_1[3] ^ (* src = "crypto_accelerator.v:4763" *) _T_2570;
  assign _T_2595 = matrix_1_1[5] ^ (* src = "crypto_accelerator.v:4764" *) matrix_1_1[2];
  assign _T_2598 = matrix_1_1[2] ^ (* src = "crypto_accelerator.v:4766" *) matrix_1_1[1];
  assign _T_2601 = matrix_1_1[5] ^ (* src = "crypto_accelerator.v:4768" *) matrix_1_1[3];
  assign _T_2604 = matrix_1_1[7] ^ (* src = "crypto_accelerator.v:4770" *) _T_2596;
  assign _T_2606 = _T_2557 ^ (* src = "crypto_accelerator.v:4771" *) _T_2596;
  assign _T_2608 = _T_2586 ^ (* src = "crypto_accelerator.v:4772" *) _T_2602;
  assign _T_2610 = _T_2562 ^ (* src = "crypto_accelerator.v:4773" *) _T_2599;
  assign _T_2612 = _T_2577 ^ (* src = "crypto_accelerator.v:4774" *) _T_2610;
  assign _T_2614 = _T_2577 ^ (* src = "crypto_accelerator.v:4775" *) _T_2599;
  assign _T_2616 = _T_2581 ^ (* src = "crypto_accelerator.v:4776" *) _T_2608;
  assign _T_2622 = _T_2614 ^ (* src = "crypto_accelerator.v:4779" *) _T_2618;
  assign _T_2626 = _T_2624 ^ (* src = "crypto_accelerator.v:4781" *) _T_2618;
  assign _T_2632 = _T_2616 ^ (* src = "crypto_accelerator.v:4784" *) _T_2628;
  assign _T_2636 = _T_2634 ^ (* src = "crypto_accelerator.v:4786" *) _T_2628;
  assign _T_2642 = _T_2640 ^ (* src = "crypto_accelerator.v:4789" *) _T_2638;
  assign _T_2646 = _T_2644 ^ (* src = "crypto_accelerator.v:4791" *) _T_2638;
  assign _T_2648 = _T_2622 ^ (* src = "crypto_accelerator.v:4792" *) _T_2620;
  assign _T_2650 = _T_2626 ^ (* src = "crypto_accelerator.v:4793" *) _T_2565;
  assign _T_2652 = _T_2632 ^ (* src = "crypto_accelerator.v:4794" *) _T_2630;
  assign _T_2654 = _T_2636 ^ (* src = "crypto_accelerator.v:4795" *) _T_2646;
  assign _T_2656 = _T_2648 ^ (* src = "crypto_accelerator.v:4796" *) _T_2642;
  assign _T_2658 = _T_2650 ^ (* src = "crypto_accelerator.v:4797" *) _T_2646;
  assign _T_2660 = _T_2652 ^ (* src = "crypto_accelerator.v:4798" *) _T_2642;
  assign _T_2662 = _T_2654 ^ (* src = "crypto_accelerator.v:4799" *) _T_2584;
  assign _T_2664 = _T_2660 ^ (* src = "crypto_accelerator.v:4800" *) _T_2662;
  assign _T_2668 = _T_2658 ^ (* src = "crypto_accelerator.v:4802" *) _T_2666;
  assign _T_2670 = _T_2656 ^ (* src = "crypto_accelerator.v:4803" *) _T_2658;
  assign _T_2672 = _T_2662 ^ (* src = "crypto_accelerator.v:4804" *) _T_2666;
  assign _T_2682 = _T_2670 ^ (* src = "crypto_accelerator.v:4809" *) _T_2666;
  assign _T_2688 = _T_2664 ^ (* src = "crypto_accelerator.v:4812" *) _T_2666;
  assign _T_2690 = _T_2658 ^ (* src = "crypto_accelerator.v:4813" *) _T_2674;
  assign _T_2692 = _T_2680 ^ (* src = "crypto_accelerator.v:4814" *) _T_2682;
  assign _T_2694 = _T_2662 ^ (* src = "crypto_accelerator.v:4815" *) _T_2676;
  assign _T_2696 = _T_2686 ^ (* src = "crypto_accelerator.v:4816" *) _T_2688;
  assign _T_2698 = _T_2692 ^ (* src = "crypto_accelerator.v:4817" *) _T_2696;
  assign _T_2700 = _T_2690 ^ (* src = "crypto_accelerator.v:4818" *) _T_2694;
  assign _T_2702 = _T_2690 ^ (* src = "crypto_accelerator.v:4819" *) _T_2692;
  assign _T_2704 = _T_2694 ^ (* src = "crypto_accelerator.v:4820" *) _T_2696;
  assign _T_2706 = _T_2700 ^ (* src = "crypto_accelerator.v:4821" *) _T_2698;
  assign _T_2744 = _T_2720 ^ (* src = "crypto_accelerator.v:4840" *) _T_2738;
  assign _T_2746 = _T_2732 ^ (* src = "crypto_accelerator.v:4841" *) _T_2734;
  assign _T_2748 = _T_2724 ^ (* src = "crypto_accelerator.v:4842" *) _T_2740;
  assign _T_2750 = _T_2710 ^ (* src = "crypto_accelerator.v:4843" *) _T_2716;
  assign _T_2752 = _T_2712 ^ (* src = "crypto_accelerator.v:4844" *) _T_2728;
  assign _T_2754 = _T_2708 ^ (* src = "crypto_accelerator.v:4845" *) _T_2718;
  assign _T_2756 = _T_2714 ^ (* src = "crypto_accelerator.v:4846" *) _T_2736;
  assign _T_2758 = _T_2744 ^ (* src = "crypto_accelerator.v:4847" *) _T_2746;
  assign _T_2760 = _T_2716 ^ (* src = "crypto_accelerator.v:4848" *) _T_2722;
  assign _T_2762 = _T_2726 ^ (* src = "crypto_accelerator.v:4849" *) _T_2742;
  assign _T_2764 = _T_2730 ^ (* src = "crypto_accelerator.v:4850" *) _T_2752;
  assign _T_2766 = _T_2744 ^ (* src = "crypto_accelerator.v:4851" *) _T_2750;
  assign _T_2768 = _T_2708 ^ (* src = "crypto_accelerator.v:4852" *) _T_2712;
  assign _T_2770 = _T_2714 ^ (* src = "crypto_accelerator.v:4853" *) _T_2718;
  assign _T_2772 = _T_2714 ^ (* src = "crypto_accelerator.v:4854" *) _T_2740;
  assign _T_2774 = _T_2724 ^ (* src = "crypto_accelerator.v:4855" *) _T_2734;
  assign _T_2776 = _T_2730 ^ (* src = "crypto_accelerator.v:4856" *) _T_2738;
  assign _T_2778 = _T_2732 ^ (* src = "crypto_accelerator.v:4857" *) _T_2748;
  assign _T_2780 = _T_2742 ^ (* src = "crypto_accelerator.v:4858" *) _T_2754;
  assign _T_2782 = _T_2748 ^ (* src = "crypto_accelerator.v:4859" *) _T_2750;
  assign _T_2784 = _T_2752 ^ (* src = "crypto_accelerator.v:4860" *) _T_2756;
  assign _T_2786 = _T_2748 ^ (* src = "crypto_accelerator.v:4861" *) _T_2758;
  assign _T_2788 = _T_2758 ^ (* src = "crypto_accelerator.v:4862" *) _T_2760;
  assign _T_2790 = _T_2754 ^ (* src = "crypto_accelerator.v:4863" *) _T_2758;
  assign _T_2792 = _T_2756 ^ (* src = "crypto_accelerator.v:4864" *) _T_2764;
  assign _T_2794 = _T_2762 ^ (* src = "crypto_accelerator.v:4865" *) _T_2766;
  assign _T_2796 = _T_2764 ^ (* src = "crypto_accelerator.v:4866" *) _T_2780;
  assign _T_2798 = _T_2766 ^ (* src = "crypto_accelerator.v:4867" *) _T_2792;
  assign _T_2800 = _T_2774 ^ (* src = "crypto_accelerator.v:4868" *) _T_2784;
  assign _T_2801 = _T_2770 ^ (* src = "crypto_accelerator.v:4869" *) _T_2786;
  assign _T_2802 = _T_2794 ^ (* src = "crypto_accelerator.v:4870" *) _T_2800;
  assign _T_2803 = _T_2778 ^ (* src = "crypto_accelerator.v:4871" *) _T_2798;
  assign _T_2804 = _T_2768 ^ (* src = "crypto_accelerator.v:4872" *) _T_2786;
  assign _T_2805 = _T_2788 ^ (* src = "crypto_accelerator.v:4873" *) _T_2796;
  assign _T_2806 = _T_2782 ^ (* src = "crypto_accelerator.v:4874" *) _T_2790;
  assign _T_2807 = _T_2772 ^ (* src = "crypto_accelerator.v:4875" *) _T_2788;
  assign _T_2808 = _T_2762 ^ (* src = "crypto_accelerator.v:4876" *) _T_2776;
  assign _T_2833 = matrix_0_2[7] ^ (* src = "crypto_accelerator.v:4878" *) matrix_0_2[4];
  assign _T_2835 = matrix_0_2[6] ^ (* src = "crypto_accelerator.v:4879" *) matrix_0_2[4];
  assign _T_2838 = matrix_0_2[7] ^ (* src = "crypto_accelerator.v:4881" *) matrix_0_2[6];
  assign _T_2841 = matrix_0_2[4] ^ (* src = "crypto_accelerator.v:4883" *) matrix_0_2[3];
  assign _T_2843 = matrix_0_2[3] ^ (* src = "crypto_accelerator.v:4884" *) matrix_0_2[0];
  assign _T_2846 = matrix_0_2[1] ^ (* src = "crypto_accelerator.v:4886" *) matrix_0_2[0];
  assign _T_2848 = matrix_0_2[6] ^ (* src = "crypto_accelerator.v:4887" *) _T_2833;
  assign _T_2851 = _T_2836 ^ (* src = "crypto_accelerator.v:4889" *) _T_2846;
  assign _T_2853 = matrix_0_2[0] ^ (* src = "crypto_accelerator.v:4890" *) _T_2841;
  assign _T_2856 = _T_2839 ^ (* src = "crypto_accelerator.v:4892" *) _T_2844;
  assign _T_2858 = _T_2839 ^ (* src = "crypto_accelerator.v:4893" *) _T_2846;
  assign _T_2860 = _T_2841 ^ (* src = "crypto_accelerator.v:4894" *) _T_2846;
  assign _T_2862 = matrix_0_2[5] ^ (* src = "crypto_accelerator.v:4895" *) _T_2841;
  assign _T_2865 = matrix_0_2[6] ^ (* src = "crypto_accelerator.v:4897" *) matrix_0_2[1];
  assign _T_2867 = matrix_0_2[5] ^ (* src = "crypto_accelerator.v:4898" *) _T_2851;
  assign _T_2870 = _T_2844 ^ (* src = "crypto_accelerator.v:4900" *) _T_2865;
  assign _T_2872 = matrix_0_2[3] ^ (* src = "crypto_accelerator.v:4901" *) _T_2849;
  assign _T_2874 = matrix_0_2[5] ^ (* src = "crypto_accelerator.v:4902" *) matrix_0_2[2];
  assign _T_2877 = matrix_0_2[2] ^ (* src = "crypto_accelerator.v:4904" *) matrix_0_2[1];
  assign _T_2880 = matrix_0_2[5] ^ (* src = "crypto_accelerator.v:4906" *) matrix_0_2[3];
  assign _T_2883 = matrix_0_2[7] ^ (* src = "crypto_accelerator.v:4908" *) _T_2875;
  assign _T_2885 = _T_2836 ^ (* src = "crypto_accelerator.v:4909" *) _T_2875;
  assign _T_2887 = _T_2865 ^ (* src = "crypto_accelerator.v:4910" *) _T_2881;
  assign _T_2889 = _T_2841 ^ (* src = "crypto_accelerator.v:4911" *) _T_2878;
  assign _T_2891 = _T_2856 ^ (* src = "crypto_accelerator.v:4912" *) _T_2889;
  assign _T_2893 = _T_2856 ^ (* src = "crypto_accelerator.v:4913" *) _T_2878;
  assign _T_2895 = _T_2860 ^ (* src = "crypto_accelerator.v:4914" *) _T_2887;
  assign _T_2901 = _T_2893 ^ (* src = "crypto_accelerator.v:4917" *) _T_2897;
  assign _T_2905 = _T_2903 ^ (* src = "crypto_accelerator.v:4919" *) _T_2897;
  assign _T_2911 = _T_2895 ^ (* src = "crypto_accelerator.v:4922" *) _T_2907;
  assign _T_2915 = _T_2913 ^ (* src = "crypto_accelerator.v:4924" *) _T_2907;
  assign _T_2921 = _T_2919 ^ (* src = "crypto_accelerator.v:4927" *) _T_2917;
  assign _T_2925 = _T_2923 ^ (* src = "crypto_accelerator.v:4929" *) _T_2917;
  assign _T_2927 = _T_2901 ^ (* src = "crypto_accelerator.v:4930" *) _T_2899;
  assign _T_2929 = _T_2905 ^ (* src = "crypto_accelerator.v:4931" *) _T_2844;
  assign _T_2931 = _T_2911 ^ (* src = "crypto_accelerator.v:4932" *) _T_2909;
  assign _T_2933 = _T_2915 ^ (* src = "crypto_accelerator.v:4933" *) _T_2925;
  assign _T_2935 = _T_2927 ^ (* src = "crypto_accelerator.v:4934" *) _T_2921;
  assign _T_2937 = _T_2929 ^ (* src = "crypto_accelerator.v:4935" *) _T_2925;
  assign _T_2939 = _T_2931 ^ (* src = "crypto_accelerator.v:4936" *) _T_2921;
  assign _T_2941 = _T_2933 ^ (* src = "crypto_accelerator.v:4937" *) _T_2863;
  assign _T_2943 = _T_2939 ^ (* src = "crypto_accelerator.v:4938" *) _T_2941;
  assign _T_2947 = _T_2937 ^ (* src = "crypto_accelerator.v:4940" *) _T_2945;
  assign _T_2949 = _T_2935 ^ (* src = "crypto_accelerator.v:4941" *) _T_2937;
  assign _T_2951 = _T_2941 ^ (* src = "crypto_accelerator.v:4942" *) _T_2945;
  assign _T_2961 = _T_2949 ^ (* src = "crypto_accelerator.v:4947" *) _T_2945;
  assign _T_2967 = _T_2943 ^ (* src = "crypto_accelerator.v:4950" *) _T_2945;
  assign _T_2969 = _T_2937 ^ (* src = "crypto_accelerator.v:4951" *) _T_2953;
  assign _T_2971 = _T_2959 ^ (* src = "crypto_accelerator.v:4952" *) _T_2961;
  assign _T_2973 = _T_2941 ^ (* src = "crypto_accelerator.v:4953" *) _T_2955;
  assign _T_2975 = _T_2965 ^ (* src = "crypto_accelerator.v:4954" *) _T_2967;
  assign _T_2977 = _T_2971 ^ (* src = "crypto_accelerator.v:4955" *) _T_2975;
  assign _T_2979 = _T_2969 ^ (* src = "crypto_accelerator.v:4956" *) _T_2973;
  assign _T_2981 = _T_2969 ^ (* src = "crypto_accelerator.v:4957" *) _T_2971;
  assign _T_2983 = _T_2973 ^ (* src = "crypto_accelerator.v:4958" *) _T_2975;
  assign _T_2985 = _T_2979 ^ (* src = "crypto_accelerator.v:4959" *) _T_2977;
  assign _T_3023 = _T_2999 ^ (* src = "crypto_accelerator.v:4978" *) _T_3017;
  assign _T_3025 = _T_3011 ^ (* src = "crypto_accelerator.v:4979" *) _T_3013;
  assign _T_3027 = _T_3003 ^ (* src = "crypto_accelerator.v:4980" *) _T_3019;
  assign _T_3029 = _T_2989 ^ (* src = "crypto_accelerator.v:4981" *) _T_2995;
  assign _T_3031 = _T_2991 ^ (* src = "crypto_accelerator.v:4982" *) _T_3007;
  assign _T_3033 = _T_2987 ^ (* src = "crypto_accelerator.v:4983" *) _T_2997;
  assign _T_3035 = _T_2993 ^ (* src = "crypto_accelerator.v:4984" *) _T_3015;
  assign _T_3037 = _T_3023 ^ (* src = "crypto_accelerator.v:4985" *) _T_3025;
  assign _T_3039 = _T_2995 ^ (* src = "crypto_accelerator.v:4986" *) _T_3001;
  assign _T_3041 = _T_3005 ^ (* src = "crypto_accelerator.v:4987" *) _T_3021;
  assign _T_3043 = _T_3009 ^ (* src = "crypto_accelerator.v:4988" *) _T_3031;
  assign _T_3045 = _T_3023 ^ (* src = "crypto_accelerator.v:4989" *) _T_3029;
  assign _T_3047 = _T_2987 ^ (* src = "crypto_accelerator.v:4990" *) _T_2991;
  assign _T_3049 = _T_2993 ^ (* src = "crypto_accelerator.v:4991" *) _T_2997;
  assign _T_3051 = _T_2993 ^ (* src = "crypto_accelerator.v:4992" *) _T_3019;
  assign _T_3053 = _T_3003 ^ (* src = "crypto_accelerator.v:4993" *) _T_3013;
  assign _T_3055 = _T_3009 ^ (* src = "crypto_accelerator.v:4994" *) _T_3017;
  assign _T_3057 = _T_3011 ^ (* src = "crypto_accelerator.v:4995" *) _T_3027;
  assign _T_3059 = _T_3021 ^ (* src = "crypto_accelerator.v:4996" *) _T_3033;
  assign _T_3061 = _T_3027 ^ (* src = "crypto_accelerator.v:4997" *) _T_3029;
  assign _T_3063 = _T_3031 ^ (* src = "crypto_accelerator.v:4998" *) _T_3035;
  assign _T_3065 = _T_3027 ^ (* src = "crypto_accelerator.v:4999" *) _T_3037;
  assign _T_3067 = _T_3037 ^ (* src = "crypto_accelerator.v:5000" *) _T_3039;
  assign _T_3069 = _T_3033 ^ (* src = "crypto_accelerator.v:5001" *) _T_3037;
  assign _T_3071 = _T_3035 ^ (* src = "crypto_accelerator.v:5002" *) _T_3043;
  assign _T_3073 = _T_3041 ^ (* src = "crypto_accelerator.v:5003" *) _T_3045;
  assign _T_3075 = _T_3043 ^ (* src = "crypto_accelerator.v:5004" *) _T_3059;
  assign _T_3077 = _T_3045 ^ (* src = "crypto_accelerator.v:5005" *) _T_3071;
  assign _T_3079 = _T_3053 ^ (* src = "crypto_accelerator.v:5006" *) _T_3063;
  assign _T_3080 = _T_3049 ^ (* src = "crypto_accelerator.v:5007" *) _T_3065;
  assign _T_3081 = _T_3073 ^ (* src = "crypto_accelerator.v:5008" *) _T_3079;
  assign _T_3082 = _T_3057 ^ (* src = "crypto_accelerator.v:5009" *) _T_3077;
  assign _T_3083 = _T_3047 ^ (* src = "crypto_accelerator.v:5010" *) _T_3065;
  assign _T_3084 = _T_3067 ^ (* src = "crypto_accelerator.v:5011" *) _T_3075;
  assign _T_3085 = _T_3061 ^ (* src = "crypto_accelerator.v:5012" *) _T_3069;
  assign _T_3086 = _T_3051 ^ (* src = "crypto_accelerator.v:5013" *) _T_3067;
  assign _T_3087 = _T_3041 ^ (* src = "crypto_accelerator.v:5014" *) _T_3055;
  assign _T_3112 = matrix_3_3[7] ^ (* src = "crypto_accelerator.v:5016" *) matrix_3_3[4];
  assign _T_3114 = matrix_3_3[6] ^ (* src = "crypto_accelerator.v:5017" *) matrix_3_3[4];
  assign _T_3117 = matrix_3_3[7] ^ (* src = "crypto_accelerator.v:5019" *) matrix_3_3[6];
  assign _T_3120 = matrix_3_3[4] ^ (* src = "crypto_accelerator.v:5021" *) matrix_3_3[3];
  assign _T_3122 = matrix_3_3[3] ^ (* src = "crypto_accelerator.v:5022" *) matrix_3_3[0];
  assign _T_3125 = matrix_3_3[1] ^ (* src = "crypto_accelerator.v:5024" *) matrix_3_3[0];
  assign _T_3127 = matrix_3_3[6] ^ (* src = "crypto_accelerator.v:5025" *) _T_3112;
  assign _T_3130 = _T_3115 ^ (* src = "crypto_accelerator.v:5027" *) _T_3125;
  assign _T_3132 = matrix_3_3[0] ^ (* src = "crypto_accelerator.v:5028" *) _T_3120;
  assign _T_3135 = _T_3118 ^ (* src = "crypto_accelerator.v:5030" *) _T_3123;
  assign _T_3137 = _T_3118 ^ (* src = "crypto_accelerator.v:5031" *) _T_3125;
  assign _T_3139 = _T_3120 ^ (* src = "crypto_accelerator.v:5032" *) _T_3125;
  assign _T_3141 = matrix_3_3[5] ^ (* src = "crypto_accelerator.v:5033" *) _T_3120;
  assign _T_3144 = matrix_3_3[6] ^ (* src = "crypto_accelerator.v:5035" *) matrix_3_3[1];
  assign _T_3146 = matrix_3_3[5] ^ (* src = "crypto_accelerator.v:5036" *) _T_3130;
  assign _T_3149 = _T_3123 ^ (* src = "crypto_accelerator.v:5038" *) _T_3144;
  assign _T_3151 = matrix_3_3[3] ^ (* src = "crypto_accelerator.v:5039" *) _T_3128;
  assign _T_3153 = matrix_3_3[5] ^ (* src = "crypto_accelerator.v:5040" *) matrix_3_3[2];
  assign _T_3156 = matrix_3_3[2] ^ (* src = "crypto_accelerator.v:5042" *) matrix_3_3[1];
  assign _T_3159 = matrix_3_3[5] ^ (* src = "crypto_accelerator.v:5044" *) matrix_3_3[3];
  assign _T_3162 = matrix_3_3[7] ^ (* src = "crypto_accelerator.v:5046" *) _T_3154;
  assign _T_3164 = _T_3115 ^ (* src = "crypto_accelerator.v:5047" *) _T_3154;
  assign _T_3166 = _T_3144 ^ (* src = "crypto_accelerator.v:5048" *) _T_3160;
  assign _T_3168 = _T_3120 ^ (* src = "crypto_accelerator.v:5049" *) _T_3157;
  assign _T_3170 = _T_3135 ^ (* src = "crypto_accelerator.v:5050" *) _T_3168;
  assign _T_3172 = _T_3135 ^ (* src = "crypto_accelerator.v:5051" *) _T_3157;
  assign _T_3174 = _T_3139 ^ (* src = "crypto_accelerator.v:5052" *) _T_3166;
  assign _T_3180 = _T_3172 ^ (* src = "crypto_accelerator.v:5055" *) _T_3176;
  assign _T_3184 = _T_3182 ^ (* src = "crypto_accelerator.v:5057" *) _T_3176;
  assign _T_3190 = _T_3174 ^ (* src = "crypto_accelerator.v:5060" *) _T_3186;
  assign _T_3194 = _T_3192 ^ (* src = "crypto_accelerator.v:5062" *) _T_3186;
  assign _T_3200 = _T_3198 ^ (* src = "crypto_accelerator.v:5065" *) _T_3196;
  assign _T_3204 = _T_3202 ^ (* src = "crypto_accelerator.v:5067" *) _T_3196;
  assign _T_3206 = _T_3180 ^ (* src = "crypto_accelerator.v:5068" *) _T_3178;
  assign _T_3208 = _T_3184 ^ (* src = "crypto_accelerator.v:5069" *) _T_3123;
  assign _T_3210 = _T_3190 ^ (* src = "crypto_accelerator.v:5070" *) _T_3188;
  assign _T_3212 = _T_3194 ^ (* src = "crypto_accelerator.v:5071" *) _T_3204;
  assign _T_3214 = _T_3206 ^ (* src = "crypto_accelerator.v:5072" *) _T_3200;
  assign _T_3216 = _T_3208 ^ (* src = "crypto_accelerator.v:5073" *) _T_3204;
  assign _T_3218 = _T_3210 ^ (* src = "crypto_accelerator.v:5074" *) _T_3200;
  assign _T_3220 = _T_3212 ^ (* src = "crypto_accelerator.v:5075" *) _T_3142;
  assign _T_3222 = _T_3218 ^ (* src = "crypto_accelerator.v:5076" *) _T_3220;
  assign _T_3226 = _T_3216 ^ (* src = "crypto_accelerator.v:5078" *) _T_3224;
  assign _T_3228 = _T_3214 ^ (* src = "crypto_accelerator.v:5079" *) _T_3216;
  assign _T_3230 = _T_3220 ^ (* src = "crypto_accelerator.v:5080" *) _T_3224;
  assign _T_3240 = _T_3228 ^ (* src = "crypto_accelerator.v:5085" *) _T_3224;
  assign _T_3246 = _T_3222 ^ (* src = "crypto_accelerator.v:5088" *) _T_3224;
  assign _T_3248 = _T_3216 ^ (* src = "crypto_accelerator.v:5089" *) _T_3232;
  assign _T_3250 = _T_3238 ^ (* src = "crypto_accelerator.v:5090" *) _T_3240;
  assign _T_3252 = _T_3220 ^ (* src = "crypto_accelerator.v:5091" *) _T_3234;
  assign _T_3254 = _T_3244 ^ (* src = "crypto_accelerator.v:5092" *) _T_3246;
  assign _T_3256 = _T_3250 ^ (* src = "crypto_accelerator.v:5093" *) _T_3254;
  assign _T_3258 = _T_3248 ^ (* src = "crypto_accelerator.v:5094" *) _T_3252;
  assign _T_3260 = _T_3248 ^ (* src = "crypto_accelerator.v:5095" *) _T_3250;
  assign _T_3262 = _T_3252 ^ (* src = "crypto_accelerator.v:5096" *) _T_3254;
  assign _T_3264 = _T_3258 ^ (* src = "crypto_accelerator.v:5097" *) _T_3256;
  assign _T_3302 = _T_3278 ^ (* src = "crypto_accelerator.v:5116" *) _T_3296;
  assign _T_3304 = _T_3290 ^ (* src = "crypto_accelerator.v:5117" *) _T_3292;
  assign _T_3306 = _T_3282 ^ (* src = "crypto_accelerator.v:5118" *) _T_3298;
  assign _T_3308 = _T_3268 ^ (* src = "crypto_accelerator.v:5119" *) _T_3274;
  assign _T_3310 = _T_3270 ^ (* src = "crypto_accelerator.v:5120" *) _T_3286;
  assign _T_3312 = _T_3266 ^ (* src = "crypto_accelerator.v:5121" *) _T_3276;
  assign _T_3314 = _T_3272 ^ (* src = "crypto_accelerator.v:5122" *) _T_3294;
  assign _T_3316 = _T_3302 ^ (* src = "crypto_accelerator.v:5123" *) _T_3304;
  assign _T_3318 = _T_3274 ^ (* src = "crypto_accelerator.v:5124" *) _T_3280;
  assign _T_3320 = _T_3284 ^ (* src = "crypto_accelerator.v:5125" *) _T_3300;
  assign _T_3322 = _T_3288 ^ (* src = "crypto_accelerator.v:5126" *) _T_3310;
  assign _T_3324 = _T_3302 ^ (* src = "crypto_accelerator.v:5127" *) _T_3308;
  assign _T_3326 = _T_3266 ^ (* src = "crypto_accelerator.v:5128" *) _T_3270;
  assign _T_3328 = _T_3272 ^ (* src = "crypto_accelerator.v:5129" *) _T_3276;
  assign _T_3330 = _T_3272 ^ (* src = "crypto_accelerator.v:5130" *) _T_3298;
  assign _T_3332 = _T_3282 ^ (* src = "crypto_accelerator.v:5131" *) _T_3292;
  assign _T_3334 = _T_3288 ^ (* src = "crypto_accelerator.v:5132" *) _T_3296;
  assign _T_3336 = _T_3290 ^ (* src = "crypto_accelerator.v:5133" *) _T_3306;
  assign _T_3338 = _T_3300 ^ (* src = "crypto_accelerator.v:5134" *) _T_3312;
  assign _T_3340 = _T_3306 ^ (* src = "crypto_accelerator.v:5135" *) _T_3308;
  assign _T_3342 = _T_3310 ^ (* src = "crypto_accelerator.v:5136" *) _T_3314;
  assign _T_3344 = _T_3306 ^ (* src = "crypto_accelerator.v:5137" *) _T_3316;
  assign _T_3346 = _T_3316 ^ (* src = "crypto_accelerator.v:5138" *) _T_3318;
  assign _T_3348 = _T_3312 ^ (* src = "crypto_accelerator.v:5139" *) _T_3316;
  assign _T_3350 = _T_3314 ^ (* src = "crypto_accelerator.v:5140" *) _T_3322;
  assign _T_3352 = _T_3320 ^ (* src = "crypto_accelerator.v:5141" *) _T_3324;
  assign _T_3354 = _T_3322 ^ (* src = "crypto_accelerator.v:5142" *) _T_3338;
  assign _T_3356 = _T_3324 ^ (* src = "crypto_accelerator.v:5143" *) _T_3350;
  assign _T_3358 = _T_3332 ^ (* src = "crypto_accelerator.v:5144" *) _T_3342;
  assign _T_3359 = _T_3328 ^ (* src = "crypto_accelerator.v:5145" *) _T_3344;
  assign _T_3360 = _T_3352 ^ (* src = "crypto_accelerator.v:5146" *) _T_3358;
  assign _T_3361 = _T_3336 ^ (* src = "crypto_accelerator.v:5147" *) _T_3356;
  assign _T_3362 = _T_3326 ^ (* src = "crypto_accelerator.v:5148" *) _T_3344;
  assign _T_3363 = _T_3346 ^ (* src = "crypto_accelerator.v:5149" *) _T_3354;
  assign _T_3364 = _T_3340 ^ (* src = "crypto_accelerator.v:5150" *) _T_3348;
  assign _T_3365 = _T_3330 ^ (* src = "crypto_accelerator.v:5151" *) _T_3346;
  assign _T_3366 = _T_3320 ^ (* src = "crypto_accelerator.v:5152" *) _T_3334;
  assign _T_3392 = matrix_3_0[7] ^ (* src = "crypto_accelerator.v:5154" *) matrix_3_0[4];
  assign _T_3394 = matrix_3_0[6] ^ (* src = "crypto_accelerator.v:5155" *) matrix_3_0[4];
  assign _T_3397 = matrix_3_0[7] ^ (* src = "crypto_accelerator.v:5157" *) matrix_3_0[6];
  assign _T_3400 = matrix_3_0[4] ^ (* src = "crypto_accelerator.v:5159" *) matrix_3_0[3];
  assign _T_3402 = matrix_3_0[3] ^ (* src = "crypto_accelerator.v:5160" *) matrix_3_0[0];
  assign _T_3405 = matrix_3_0[1] ^ (* src = "crypto_accelerator.v:5162" *) matrix_3_0[0];
  assign _T_3407 = matrix_3_0[6] ^ (* src = "crypto_accelerator.v:5163" *) _T_3392;
  assign _T_3410 = _T_3395 ^ (* src = "crypto_accelerator.v:5165" *) _T_3405;
  assign _T_3412 = matrix_3_0[0] ^ (* src = "crypto_accelerator.v:5166" *) _T_3400;
  assign _T_3415 = _T_3398 ^ (* src = "crypto_accelerator.v:5168" *) _T_3403;
  assign _T_3417 = _T_3398 ^ (* src = "crypto_accelerator.v:5169" *) _T_3405;
  assign _T_3419 = _T_3400 ^ (* src = "crypto_accelerator.v:5170" *) _T_3405;
  assign _T_3421 = matrix_3_0[5] ^ (* src = "crypto_accelerator.v:5171" *) _T_3400;
  assign _T_3424 = matrix_3_0[6] ^ (* src = "crypto_accelerator.v:5173" *) matrix_3_0[1];
  assign _T_3426 = matrix_3_0[5] ^ (* src = "crypto_accelerator.v:5174" *) _T_3410;
  assign _T_3429 = _T_3403 ^ (* src = "crypto_accelerator.v:5176" *) _T_3424;
  assign _T_3431 = matrix_3_0[3] ^ (* src = "crypto_accelerator.v:5177" *) _T_3408;
  assign _T_3433 = matrix_3_0[5] ^ (* src = "crypto_accelerator.v:5178" *) matrix_3_0[2];
  assign _T_3436 = matrix_3_0[2] ^ (* src = "crypto_accelerator.v:5180" *) matrix_3_0[1];
  assign _T_3439 = matrix_3_0[5] ^ (* src = "crypto_accelerator.v:5182" *) matrix_3_0[3];
  assign _T_3442 = matrix_3_0[7] ^ (* src = "crypto_accelerator.v:5184" *) _T_3434;
  assign _T_3444 = _T_3395 ^ (* src = "crypto_accelerator.v:5185" *) _T_3434;
  assign _T_3446 = _T_3424 ^ (* src = "crypto_accelerator.v:5186" *) _T_3440;
  assign _T_3448 = _T_3400 ^ (* src = "crypto_accelerator.v:5187" *) _T_3437;
  assign _T_3450 = _T_3415 ^ (* src = "crypto_accelerator.v:5188" *) _T_3448;
  assign _T_3452 = _T_3415 ^ (* src = "crypto_accelerator.v:5189" *) _T_3437;
  assign _T_3454 = _T_3419 ^ (* src = "crypto_accelerator.v:5190" *) _T_3446;
  assign _T_3460 = _T_3452 ^ (* src = "crypto_accelerator.v:5193" *) _T_3456;
  assign _T_3464 = _T_3462 ^ (* src = "crypto_accelerator.v:5195" *) _T_3456;
  assign _T_3470 = _T_3454 ^ (* src = "crypto_accelerator.v:5198" *) _T_3466;
  assign _T_3474 = _T_3472 ^ (* src = "crypto_accelerator.v:5200" *) _T_3466;
  assign _T_3480 = _T_3478 ^ (* src = "crypto_accelerator.v:5203" *) _T_3476;
  assign _T_3484 = _T_3482 ^ (* src = "crypto_accelerator.v:5205" *) _T_3476;
  assign _T_3486 = _T_3460 ^ (* src = "crypto_accelerator.v:5206" *) _T_3458;
  assign _T_3488 = _T_3464 ^ (* src = "crypto_accelerator.v:5207" *) _T_3403;
  assign _T_3490 = _T_3470 ^ (* src = "crypto_accelerator.v:5208" *) _T_3468;
  assign _T_3492 = _T_3474 ^ (* src = "crypto_accelerator.v:5209" *) _T_3484;
  assign _T_3494 = _T_3486 ^ (* src = "crypto_accelerator.v:5210" *) _T_3480;
  assign _T_3496 = _T_3488 ^ (* src = "crypto_accelerator.v:5211" *) _T_3484;
  assign _T_3498 = _T_3490 ^ (* src = "crypto_accelerator.v:5212" *) _T_3480;
  assign _T_3500 = _T_3492 ^ (* src = "crypto_accelerator.v:5213" *) _T_3422;
  assign _T_3502 = _T_3498 ^ (* src = "crypto_accelerator.v:5214" *) _T_3500;
  assign _T_3506 = _T_3496 ^ (* src = "crypto_accelerator.v:5216" *) _T_3504;
  assign _T_3508 = _T_3494 ^ (* src = "crypto_accelerator.v:5217" *) _T_3496;
  assign _T_3510 = _T_3500 ^ (* src = "crypto_accelerator.v:5218" *) _T_3504;
  assign _T_3520 = _T_3508 ^ (* src = "crypto_accelerator.v:5223" *) _T_3504;
  assign _T_3526 = _T_3502 ^ (* src = "crypto_accelerator.v:5226" *) _T_3504;
  assign _T_3528 = _T_3496 ^ (* src = "crypto_accelerator.v:5227" *) _T_3512;
  assign _T_3530 = _T_3518 ^ (* src = "crypto_accelerator.v:5228" *) _T_3520;
  assign _T_3532 = _T_3500 ^ (* src = "crypto_accelerator.v:5229" *) _T_3514;
  assign _T_3534 = _T_3524 ^ (* src = "crypto_accelerator.v:5230" *) _T_3526;
  assign _T_3536 = _T_3530 ^ (* src = "crypto_accelerator.v:5231" *) _T_3534;
  assign _T_3538 = _T_3528 ^ (* src = "crypto_accelerator.v:5232" *) _T_3532;
  assign _T_3540 = _T_3528 ^ (* src = "crypto_accelerator.v:5233" *) _T_3530;
  assign _T_3542 = _T_3532 ^ (* src = "crypto_accelerator.v:5234" *) _T_3534;
  assign _T_3544 = _T_3538 ^ (* src = "crypto_accelerator.v:5235" *) _T_3536;
  assign _T_3582 = _T_3558 ^ (* src = "crypto_accelerator.v:5254" *) _T_3576;
  assign _T_3584 = _T_3570 ^ (* src = "crypto_accelerator.v:5255" *) _T_3572;
  assign _T_3586 = _T_3562 ^ (* src = "crypto_accelerator.v:5256" *) _T_3578;
  assign _T_3588 = _T_3548 ^ (* src = "crypto_accelerator.v:5257" *) _T_3554;
  assign _T_3590 = _T_3550 ^ (* src = "crypto_accelerator.v:5258" *) _T_3566;
  assign _T_3592 = _T_3546 ^ (* src = "crypto_accelerator.v:5259" *) _T_3556;
  assign _T_3594 = _T_3552 ^ (* src = "crypto_accelerator.v:5260" *) _T_3574;
  assign _T_3596 = _T_3582 ^ (* src = "crypto_accelerator.v:5261" *) _T_3584;
  assign _T_3598 = _T_3554 ^ (* src = "crypto_accelerator.v:5262" *) _T_3560;
  assign _T_3600 = _T_3564 ^ (* src = "crypto_accelerator.v:5263" *) _T_3580;
  assign _T_3602 = _T_3568 ^ (* src = "crypto_accelerator.v:5264" *) _T_3590;
  assign _T_3604 = _T_3582 ^ (* src = "crypto_accelerator.v:5265" *) _T_3588;
  assign _T_3606 = _T_3546 ^ (* src = "crypto_accelerator.v:5266" *) _T_3550;
  assign _T_3608 = _T_3552 ^ (* src = "crypto_accelerator.v:5267" *) _T_3556;
  assign _T_3610 = _T_3552 ^ (* src = "crypto_accelerator.v:5268" *) _T_3578;
  assign _T_3612 = _T_3562 ^ (* src = "crypto_accelerator.v:5269" *) _T_3572;
  assign _T_3614 = _T_3568 ^ (* src = "crypto_accelerator.v:5270" *) _T_3576;
  assign _T_3616 = _T_3570 ^ (* src = "crypto_accelerator.v:5271" *) _T_3586;
  assign _T_3618 = _T_3580 ^ (* src = "crypto_accelerator.v:5272" *) _T_3592;
  assign _T_3620 = _T_3586 ^ (* src = "crypto_accelerator.v:5273" *) _T_3588;
  assign _T_3622 = _T_3590 ^ (* src = "crypto_accelerator.v:5274" *) _T_3594;
  assign _T_3624 = _T_3586 ^ (* src = "crypto_accelerator.v:5275" *) _T_3596;
  assign _T_3626 = _T_3596 ^ (* src = "crypto_accelerator.v:5276" *) _T_3598;
  assign _T_3628 = _T_3592 ^ (* src = "crypto_accelerator.v:5277" *) _T_3596;
  assign _T_3630 = _T_3594 ^ (* src = "crypto_accelerator.v:5278" *) _T_3602;
  assign _T_3632 = _T_3600 ^ (* src = "crypto_accelerator.v:5279" *) _T_3604;
  assign _T_3634 = _T_3602 ^ (* src = "crypto_accelerator.v:5280" *) _T_3618;
  assign _T_3636 = _T_3604 ^ (* src = "crypto_accelerator.v:5281" *) _T_3630;
  assign _T_3638 = _T_3612 ^ (* src = "crypto_accelerator.v:5282" *) _T_3622;
  assign _T_3639 = _T_3608 ^ (* src = "crypto_accelerator.v:5283" *) _T_3624;
  assign _T_3640 = _T_3632 ^ (* src = "crypto_accelerator.v:5284" *) _T_3638;
  assign _T_3641 = _T_3616 ^ (* src = "crypto_accelerator.v:5285" *) _T_3636;
  assign _T_3642 = _T_3606 ^ (* src = "crypto_accelerator.v:5286" *) _T_3624;
  assign _T_3643 = _T_3626 ^ (* src = "crypto_accelerator.v:5287" *) _T_3634;
  assign _T_3644 = _T_3620 ^ (* src = "crypto_accelerator.v:5288" *) _T_3628;
  assign _T_3645 = _T_3610 ^ (* src = "crypto_accelerator.v:5289" *) _T_3626;
  assign _T_3646 = _T_3600 ^ (* src = "crypto_accelerator.v:5290" *) _T_3614;
  assign _T_3671 = matrix_2_1[7] ^ (* src = "crypto_accelerator.v:5292" *) matrix_2_1[4];
  assign _T_3673 = matrix_2_1[6] ^ (* src = "crypto_accelerator.v:5293" *) matrix_2_1[4];
  assign _T_3676 = matrix_2_1[7] ^ (* src = "crypto_accelerator.v:5295" *) matrix_2_1[6];
  assign _T_3679 = matrix_2_1[4] ^ (* src = "crypto_accelerator.v:5297" *) matrix_2_1[3];
  assign _T_3681 = matrix_2_1[3] ^ (* src = "crypto_accelerator.v:5298" *) matrix_2_1[0];
  assign _T_3684 = matrix_2_1[1] ^ (* src = "crypto_accelerator.v:5300" *) matrix_2_1[0];
  assign _T_3686 = matrix_2_1[6] ^ (* src = "crypto_accelerator.v:5301" *) _T_3671;
  assign _T_3689 = _T_3674 ^ (* src = "crypto_accelerator.v:5303" *) _T_3684;
  assign _T_3691 = matrix_2_1[0] ^ (* src = "crypto_accelerator.v:5304" *) _T_3679;
  assign _T_3694 = _T_3677 ^ (* src = "crypto_accelerator.v:5306" *) _T_3682;
  assign _T_3696 = _T_3677 ^ (* src = "crypto_accelerator.v:5307" *) _T_3684;
  assign _T_3698 = _T_3679 ^ (* src = "crypto_accelerator.v:5308" *) _T_3684;
  assign _T_3700 = matrix_2_1[5] ^ (* src = "crypto_accelerator.v:5309" *) _T_3679;
  assign _T_3703 = matrix_2_1[6] ^ (* src = "crypto_accelerator.v:5311" *) matrix_2_1[1];
  assign _T_3705 = matrix_2_1[5] ^ (* src = "crypto_accelerator.v:5312" *) _T_3689;
  assign _T_3708 = _T_3682 ^ (* src = "crypto_accelerator.v:5314" *) _T_3703;
  assign _T_3710 = matrix_2_1[3] ^ (* src = "crypto_accelerator.v:5315" *) _T_3687;
  assign _T_3712 = matrix_2_1[5] ^ (* src = "crypto_accelerator.v:5316" *) matrix_2_1[2];
  assign _T_3715 = matrix_2_1[2] ^ (* src = "crypto_accelerator.v:5318" *) matrix_2_1[1];
  assign _T_3718 = matrix_2_1[5] ^ (* src = "crypto_accelerator.v:5320" *) matrix_2_1[3];
  assign _T_3721 = matrix_2_1[7] ^ (* src = "crypto_accelerator.v:5322" *) _T_3713;
  assign _T_3723 = _T_3674 ^ (* src = "crypto_accelerator.v:5323" *) _T_3713;
  assign _T_3725 = _T_3703 ^ (* src = "crypto_accelerator.v:5324" *) _T_3719;
  assign _T_3727 = _T_3679 ^ (* src = "crypto_accelerator.v:5325" *) _T_3716;
  assign _T_3729 = _T_3694 ^ (* src = "crypto_accelerator.v:5326" *) _T_3727;
  assign _T_3731 = _T_3694 ^ (* src = "crypto_accelerator.v:5327" *) _T_3716;
  assign _T_3733 = _T_3698 ^ (* src = "crypto_accelerator.v:5328" *) _T_3725;
  assign _T_3739 = _T_3731 ^ (* src = "crypto_accelerator.v:5331" *) _T_3735;
  assign _T_3743 = _T_3741 ^ (* src = "crypto_accelerator.v:5333" *) _T_3735;
  assign _T_3749 = _T_3733 ^ (* src = "crypto_accelerator.v:5336" *) _T_3745;
  assign _T_3753 = _T_3751 ^ (* src = "crypto_accelerator.v:5338" *) _T_3745;
  assign _T_3759 = _T_3757 ^ (* src = "crypto_accelerator.v:5341" *) _T_3755;
  assign _T_3763 = _T_3761 ^ (* src = "crypto_accelerator.v:5343" *) _T_3755;
  assign _T_3765 = _T_3739 ^ (* src = "crypto_accelerator.v:5344" *) _T_3737;
  assign _T_3767 = _T_3743 ^ (* src = "crypto_accelerator.v:5345" *) _T_3682;
  assign _T_3769 = _T_3749 ^ (* src = "crypto_accelerator.v:5346" *) _T_3747;
  assign _T_3771 = _T_3753 ^ (* src = "crypto_accelerator.v:5347" *) _T_3763;
  assign _T_3773 = _T_3765 ^ (* src = "crypto_accelerator.v:5348" *) _T_3759;
  assign _T_3775 = _T_3767 ^ (* src = "crypto_accelerator.v:5349" *) _T_3763;
  assign _T_3777 = _T_3769 ^ (* src = "crypto_accelerator.v:5350" *) _T_3759;
  assign _T_3779 = _T_3771 ^ (* src = "crypto_accelerator.v:5351" *) _T_3701;
  assign _T_3781 = _T_3777 ^ (* src = "crypto_accelerator.v:5352" *) _T_3779;
  assign _T_3785 = _T_3775 ^ (* src = "crypto_accelerator.v:5354" *) _T_3783;
  assign _T_3787 = _T_3773 ^ (* src = "crypto_accelerator.v:5355" *) _T_3775;
  assign _T_3789 = _T_3779 ^ (* src = "crypto_accelerator.v:5356" *) _T_3783;
  assign _T_3799 = _T_3787 ^ (* src = "crypto_accelerator.v:5361" *) _T_3783;
  assign _T_3805 = _T_3781 ^ (* src = "crypto_accelerator.v:5364" *) _T_3783;
  assign _T_3807 = _T_3775 ^ (* src = "crypto_accelerator.v:5365" *) _T_3791;
  assign _T_3809 = _T_3797 ^ (* src = "crypto_accelerator.v:5366" *) _T_3799;
  assign _T_3811 = _T_3779 ^ (* src = "crypto_accelerator.v:5367" *) _T_3793;
  assign _T_3813 = _T_3803 ^ (* src = "crypto_accelerator.v:5368" *) _T_3805;
  assign _T_3815 = _T_3809 ^ (* src = "crypto_accelerator.v:5369" *) _T_3813;
  assign _T_3817 = _T_3807 ^ (* src = "crypto_accelerator.v:5370" *) _T_3811;
  assign _T_3819 = _T_3807 ^ (* src = "crypto_accelerator.v:5371" *) _T_3809;
  assign _T_3821 = _T_3811 ^ (* src = "crypto_accelerator.v:5372" *) _T_3813;
  assign _T_3823 = _T_3817 ^ (* src = "crypto_accelerator.v:5373" *) _T_3815;
  assign _T_3861 = _T_3837 ^ (* src = "crypto_accelerator.v:5392" *) _T_3855;
  assign _T_3863 = _T_3849 ^ (* src = "crypto_accelerator.v:5393" *) _T_3851;
  assign _T_3865 = _T_3841 ^ (* src = "crypto_accelerator.v:5394" *) _T_3857;
  assign _T_3867 = _T_3827 ^ (* src = "crypto_accelerator.v:5395" *) _T_3833;
  assign _T_3869 = _T_3829 ^ (* src = "crypto_accelerator.v:5396" *) _T_3845;
  assign _T_3871 = _T_3825 ^ (* src = "crypto_accelerator.v:5397" *) _T_3835;
  assign _T_3873 = _T_3831 ^ (* src = "crypto_accelerator.v:5398" *) _T_3853;
  assign _T_3875 = _T_3861 ^ (* src = "crypto_accelerator.v:5399" *) _T_3863;
  assign _T_3877 = _T_3833 ^ (* src = "crypto_accelerator.v:5400" *) _T_3839;
  assign _T_3879 = _T_3843 ^ (* src = "crypto_accelerator.v:5401" *) _T_3859;
  assign _T_3881 = _T_3847 ^ (* src = "crypto_accelerator.v:5402" *) _T_3869;
  assign _T_3883 = _T_3861 ^ (* src = "crypto_accelerator.v:5403" *) _T_3867;
  assign _T_3885 = _T_3825 ^ (* src = "crypto_accelerator.v:5404" *) _T_3829;
  assign _T_3887 = _T_3831 ^ (* src = "crypto_accelerator.v:5405" *) _T_3835;
  assign _T_3889 = _T_3831 ^ (* src = "crypto_accelerator.v:5406" *) _T_3857;
  assign _T_3891 = _T_3841 ^ (* src = "crypto_accelerator.v:5407" *) _T_3851;
  assign _T_3893 = _T_3847 ^ (* src = "crypto_accelerator.v:5408" *) _T_3855;
  assign _T_3895 = _T_3849 ^ (* src = "crypto_accelerator.v:5409" *) _T_3865;
  assign _T_3897 = _T_3859 ^ (* src = "crypto_accelerator.v:5410" *) _T_3871;
  assign _T_3899 = _T_3865 ^ (* src = "crypto_accelerator.v:5411" *) _T_3867;
  assign _T_3901 = _T_3869 ^ (* src = "crypto_accelerator.v:5412" *) _T_3873;
  assign _T_3903 = _T_3865 ^ (* src = "crypto_accelerator.v:5413" *) _T_3875;
  assign _T_3905 = _T_3875 ^ (* src = "crypto_accelerator.v:5414" *) _T_3877;
  assign _T_3907 = _T_3871 ^ (* src = "crypto_accelerator.v:5415" *) _T_3875;
  assign _T_3909 = _T_3873 ^ (* src = "crypto_accelerator.v:5416" *) _T_3881;
  assign _T_3911 = _T_3879 ^ (* src = "crypto_accelerator.v:5417" *) _T_3883;
  assign _T_3913 = _T_3881 ^ (* src = "crypto_accelerator.v:5418" *) _T_3897;
  assign _T_3915 = _T_3883 ^ (* src = "crypto_accelerator.v:5419" *) _T_3909;
  assign _T_3917 = _T_3891 ^ (* src = "crypto_accelerator.v:5420" *) _T_3901;
  assign _T_3918 = _T_3887 ^ (* src = "crypto_accelerator.v:5421" *) _T_3903;
  assign _T_3919 = _T_3911 ^ (* src = "crypto_accelerator.v:5422" *) _T_3917;
  assign _T_3920 = _T_3895 ^ (* src = "crypto_accelerator.v:5423" *) _T_3915;
  assign _T_3921 = _T_3885 ^ (* src = "crypto_accelerator.v:5424" *) _T_3903;
  assign _T_3922 = _T_3905 ^ (* src = "crypto_accelerator.v:5425" *) _T_3913;
  assign _T_3923 = _T_3899 ^ (* src = "crypto_accelerator.v:5426" *) _T_3907;
  assign _T_3924 = _T_3889 ^ (* src = "crypto_accelerator.v:5427" *) _T_3905;
  assign _T_3925 = _T_3879 ^ (* src = "crypto_accelerator.v:5428" *) _T_3893;
  assign _T_3950 = matrix_1_2[7] ^ (* src = "crypto_accelerator.v:5430" *) matrix_1_2[4];
  assign _T_3952 = matrix_1_2[6] ^ (* src = "crypto_accelerator.v:5431" *) matrix_1_2[4];
  assign _T_3955 = matrix_1_2[7] ^ (* src = "crypto_accelerator.v:5433" *) matrix_1_2[6];
  assign _T_3958 = matrix_1_2[4] ^ (* src = "crypto_accelerator.v:5435" *) matrix_1_2[3];
  assign _T_3960 = matrix_1_2[3] ^ (* src = "crypto_accelerator.v:5436" *) matrix_1_2[0];
  assign _T_3963 = matrix_1_2[1] ^ (* src = "crypto_accelerator.v:5438" *) matrix_1_2[0];
  assign _T_3965 = matrix_1_2[6] ^ (* src = "crypto_accelerator.v:5439" *) _T_3950;
  assign _T_3968 = _T_3953 ^ (* src = "crypto_accelerator.v:5441" *) _T_3963;
  assign _T_3970 = matrix_1_2[0] ^ (* src = "crypto_accelerator.v:5442" *) _T_3958;
  assign _T_3973 = _T_3956 ^ (* src = "crypto_accelerator.v:5444" *) _T_3961;
  assign _T_3975 = _T_3956 ^ (* src = "crypto_accelerator.v:5445" *) _T_3963;
  assign _T_3977 = _T_3958 ^ (* src = "crypto_accelerator.v:5446" *) _T_3963;
  assign _T_3979 = matrix_1_2[5] ^ (* src = "crypto_accelerator.v:5447" *) _T_3958;
  assign _T_3982 = matrix_1_2[6] ^ (* src = "crypto_accelerator.v:5449" *) matrix_1_2[1];
  assign _T_3984 = matrix_1_2[5] ^ (* src = "crypto_accelerator.v:5450" *) _T_3968;
  assign _T_3987 = _T_3961 ^ (* src = "crypto_accelerator.v:5452" *) _T_3982;
  assign _T_3989 = matrix_1_2[3] ^ (* src = "crypto_accelerator.v:5453" *) _T_3966;
  assign _T_3991 = matrix_1_2[5] ^ (* src = "crypto_accelerator.v:5454" *) matrix_1_2[2];
  assign _T_3994 = matrix_1_2[2] ^ (* src = "crypto_accelerator.v:5456" *) matrix_1_2[1];
  assign _T_3997 = matrix_1_2[5] ^ (* src = "crypto_accelerator.v:5458" *) matrix_1_2[3];
  assign _T_4000 = matrix_1_2[7] ^ (* src = "crypto_accelerator.v:5460" *) _T_3992;
  assign _T_4002 = _T_3953 ^ (* src = "crypto_accelerator.v:5461" *) _T_3992;
  assign _T_4004 = _T_3982 ^ (* src = "crypto_accelerator.v:5462" *) _T_3998;
  assign _T_4006 = _T_3958 ^ (* src = "crypto_accelerator.v:5463" *) _T_3995;
  assign _T_4008 = _T_3973 ^ (* src = "crypto_accelerator.v:5464" *) _T_4006;
  assign _T_4010 = _T_3973 ^ (* src = "crypto_accelerator.v:5465" *) _T_3995;
  assign _T_4012 = _T_3977 ^ (* src = "crypto_accelerator.v:5466" *) _T_4004;
  assign _T_4018 = _T_4010 ^ (* src = "crypto_accelerator.v:5469" *) _T_4014;
  assign _T_4022 = _T_4020 ^ (* src = "crypto_accelerator.v:5471" *) _T_4014;
  assign _T_4028 = _T_4012 ^ (* src = "crypto_accelerator.v:5474" *) _T_4024;
  assign _T_4032 = _T_4030 ^ (* src = "crypto_accelerator.v:5476" *) _T_4024;
  assign _T_4038 = _T_4036 ^ (* src = "crypto_accelerator.v:5479" *) _T_4034;
  assign _T_4042 = _T_4040 ^ (* src = "crypto_accelerator.v:5481" *) _T_4034;
  assign _T_4044 = _T_4018 ^ (* src = "crypto_accelerator.v:5482" *) _T_4016;
  assign _T_4046 = _T_4022 ^ (* src = "crypto_accelerator.v:5483" *) _T_3961;
  assign _T_4048 = _T_4028 ^ (* src = "crypto_accelerator.v:5484" *) _T_4026;
  assign _T_4050 = _T_4032 ^ (* src = "crypto_accelerator.v:5485" *) _T_4042;
  assign _T_4052 = _T_4044 ^ (* src = "crypto_accelerator.v:5486" *) _T_4038;
  assign _T_4054 = _T_4046 ^ (* src = "crypto_accelerator.v:5487" *) _T_4042;
  assign _T_4056 = _T_4048 ^ (* src = "crypto_accelerator.v:5488" *) _T_4038;
  assign _T_4058 = _T_4050 ^ (* src = "crypto_accelerator.v:5489" *) _T_3980;
  assign _T_4060 = _T_4056 ^ (* src = "crypto_accelerator.v:5490" *) _T_4058;
  assign _T_4064 = _T_4054 ^ (* src = "crypto_accelerator.v:5492" *) _T_4062;
  assign _T_4066 = _T_4052 ^ (* src = "crypto_accelerator.v:5493" *) _T_4054;
  assign _T_4068 = _T_4058 ^ (* src = "crypto_accelerator.v:5494" *) _T_4062;
  assign _T_4078 = _T_4066 ^ (* src = "crypto_accelerator.v:5499" *) _T_4062;
  assign _T_4084 = _T_4060 ^ (* src = "crypto_accelerator.v:5502" *) _T_4062;
  assign _T_4086 = _T_4054 ^ (* src = "crypto_accelerator.v:5503" *) _T_4070;
  assign _T_4088 = _T_4076 ^ (* src = "crypto_accelerator.v:5504" *) _T_4078;
  assign _T_4090 = _T_4058 ^ (* src = "crypto_accelerator.v:5505" *) _T_4072;
  assign _T_4092 = _T_4082 ^ (* src = "crypto_accelerator.v:5506" *) _T_4084;
  assign _T_4094 = _T_4088 ^ (* src = "crypto_accelerator.v:5507" *) _T_4092;
  assign _T_4096 = _T_4086 ^ (* src = "crypto_accelerator.v:5508" *) _T_4090;
  assign _T_4098 = _T_4086 ^ (* src = "crypto_accelerator.v:5509" *) _T_4088;
  assign _T_4100 = _T_4090 ^ (* src = "crypto_accelerator.v:5510" *) _T_4092;
  assign _T_4102 = _T_4096 ^ (* src = "crypto_accelerator.v:5511" *) _T_4094;
  assign _T_4140 = _T_4116 ^ (* src = "crypto_accelerator.v:5530" *) _T_4134;
  assign _T_4142 = _T_4128 ^ (* src = "crypto_accelerator.v:5531" *) _T_4130;
  assign _T_4144 = _T_4120 ^ (* src = "crypto_accelerator.v:5532" *) _T_4136;
  assign _T_4146 = _T_4106 ^ (* src = "crypto_accelerator.v:5533" *) _T_4112;
  assign _T_4148 = _T_4108 ^ (* src = "crypto_accelerator.v:5534" *) _T_4124;
  assign _T_4150 = _T_4104 ^ (* src = "crypto_accelerator.v:5535" *) _T_4114;
  assign _T_4152 = _T_4110 ^ (* src = "crypto_accelerator.v:5536" *) _T_4132;
  assign _T_4154 = _T_4140 ^ (* src = "crypto_accelerator.v:5537" *) _T_4142;
  assign _T_4156 = _T_4112 ^ (* src = "crypto_accelerator.v:5538" *) _T_4118;
  assign _T_4158 = _T_4122 ^ (* src = "crypto_accelerator.v:5539" *) _T_4138;
  assign _T_4160 = _T_4126 ^ (* src = "crypto_accelerator.v:5540" *) _T_4148;
  assign _T_4162 = _T_4140 ^ (* src = "crypto_accelerator.v:5541" *) _T_4146;
  assign _T_4164 = _T_4104 ^ (* src = "crypto_accelerator.v:5542" *) _T_4108;
  assign _T_4166 = _T_4110 ^ (* src = "crypto_accelerator.v:5543" *) _T_4114;
  assign _T_4168 = _T_4110 ^ (* src = "crypto_accelerator.v:5544" *) _T_4136;
  assign _T_4170 = _T_4120 ^ (* src = "crypto_accelerator.v:5545" *) _T_4130;
  assign _T_4172 = _T_4126 ^ (* src = "crypto_accelerator.v:5546" *) _T_4134;
  assign _T_4174 = _T_4128 ^ (* src = "crypto_accelerator.v:5547" *) _T_4144;
  assign _T_4176 = _T_4138 ^ (* src = "crypto_accelerator.v:5548" *) _T_4150;
  assign _T_4178 = _T_4144 ^ (* src = "crypto_accelerator.v:5549" *) _T_4146;
  assign _T_4180 = _T_4148 ^ (* src = "crypto_accelerator.v:5550" *) _T_4152;
  assign _T_4182 = _T_4144 ^ (* src = "crypto_accelerator.v:5551" *) _T_4154;
  assign _T_4184 = _T_4154 ^ (* src = "crypto_accelerator.v:5552" *) _T_4156;
  assign _T_4186 = _T_4150 ^ (* src = "crypto_accelerator.v:5553" *) _T_4154;
  assign _T_4188 = _T_4152 ^ (* src = "crypto_accelerator.v:5554" *) _T_4160;
  assign _T_4190 = _T_4158 ^ (* src = "crypto_accelerator.v:5555" *) _T_4162;
  assign _T_4192 = _T_4160 ^ (* src = "crypto_accelerator.v:5556" *) _T_4176;
  assign _T_4194 = _T_4162 ^ (* src = "crypto_accelerator.v:5557" *) _T_4188;
  assign _T_4196 = _T_4170 ^ (* src = "crypto_accelerator.v:5558" *) _T_4180;
  assign _T_4197 = _T_4166 ^ (* src = "crypto_accelerator.v:5559" *) _T_4182;
  assign _T_4198 = _T_4190 ^ (* src = "crypto_accelerator.v:5560" *) _T_4196;
  assign _T_4199 = _T_4174 ^ (* src = "crypto_accelerator.v:5561" *) _T_4194;
  assign _T_4200 = _T_4164 ^ (* src = "crypto_accelerator.v:5562" *) _T_4182;
  assign _T_4201 = _T_4184 ^ (* src = "crypto_accelerator.v:5563" *) _T_4192;
  assign _T_4202 = _T_4178 ^ (* src = "crypto_accelerator.v:5564" *) _T_4186;
  assign _T_4203 = _T_4168 ^ (* src = "crypto_accelerator.v:5565" *) _T_4184;
  assign _T_4204 = _T_4158 ^ (* src = "crypto_accelerator.v:5566" *) _T_4172;
  assign _T_4229 = matrix_0_3[7] ^ (* src = "crypto_accelerator.v:5568" *) matrix_0_3[4];
  assign _T_4231 = matrix_0_3[6] ^ (* src = "crypto_accelerator.v:5569" *) matrix_0_3[4];
  assign _T_4234 = matrix_0_3[7] ^ (* src = "crypto_accelerator.v:5571" *) matrix_0_3[6];
  assign _T_4237 = matrix_0_3[4] ^ (* src = "crypto_accelerator.v:5573" *) matrix_0_3[3];
  assign _T_4239 = matrix_0_3[3] ^ (* src = "crypto_accelerator.v:5574" *) matrix_0_3[0];
  assign _T_4242 = matrix_0_3[1] ^ (* src = "crypto_accelerator.v:5576" *) matrix_0_3[0];
  assign _T_4244 = matrix_0_3[6] ^ (* src = "crypto_accelerator.v:5577" *) _T_4229;
  assign _T_4247 = _T_4232 ^ (* src = "crypto_accelerator.v:5579" *) _T_4242;
  assign _T_4249 = matrix_0_3[0] ^ (* src = "crypto_accelerator.v:5580" *) _T_4237;
  assign _T_4252 = _T_4235 ^ (* src = "crypto_accelerator.v:5582" *) _T_4240;
  assign _T_4254 = _T_4235 ^ (* src = "crypto_accelerator.v:5583" *) _T_4242;
  assign _T_4256 = _T_4237 ^ (* src = "crypto_accelerator.v:5584" *) _T_4242;
  assign _T_4258 = matrix_0_3[5] ^ (* src = "crypto_accelerator.v:5585" *) _T_4237;
  assign _T_4261 = matrix_0_3[6] ^ (* src = "crypto_accelerator.v:5587" *) matrix_0_3[1];
  assign _T_4263 = matrix_0_3[5] ^ (* src = "crypto_accelerator.v:5588" *) _T_4247;
  assign _T_4266 = _T_4240 ^ (* src = "crypto_accelerator.v:5590" *) _T_4261;
  assign _T_4268 = matrix_0_3[3] ^ (* src = "crypto_accelerator.v:5591" *) _T_4245;
  assign _T_4270 = matrix_0_3[5] ^ (* src = "crypto_accelerator.v:5592" *) matrix_0_3[2];
  assign _T_4273 = matrix_0_3[2] ^ (* src = "crypto_accelerator.v:5594" *) matrix_0_3[1];
  assign _T_4276 = matrix_0_3[5] ^ (* src = "crypto_accelerator.v:5596" *) matrix_0_3[3];
  assign _T_4279 = matrix_0_3[7] ^ (* src = "crypto_accelerator.v:5598" *) _T_4271;
  assign _T_4281 = _T_4232 ^ (* src = "crypto_accelerator.v:5599" *) _T_4271;
  assign _T_4283 = _T_4261 ^ (* src = "crypto_accelerator.v:5600" *) _T_4277;
  assign _T_4285 = _T_4237 ^ (* src = "crypto_accelerator.v:5601" *) _T_4274;
  assign _T_4287 = _T_4252 ^ (* src = "crypto_accelerator.v:5602" *) _T_4285;
  assign _T_4289 = _T_4252 ^ (* src = "crypto_accelerator.v:5603" *) _T_4274;
  assign _T_4291 = _T_4256 ^ (* src = "crypto_accelerator.v:5604" *) _T_4283;
  assign _T_4297 = _T_4289 ^ (* src = "crypto_accelerator.v:5607" *) _T_4293;
  assign _T_4301 = _T_4299 ^ (* src = "crypto_accelerator.v:5609" *) _T_4293;
  assign _T_4307 = _T_4291 ^ (* src = "crypto_accelerator.v:5612" *) _T_4303;
  assign _T_4311 = _T_4309 ^ (* src = "crypto_accelerator.v:5614" *) _T_4303;
  assign _T_4317 = _T_4315 ^ (* src = "crypto_accelerator.v:5617" *) _T_4313;
  assign _T_4321 = _T_4319 ^ (* src = "crypto_accelerator.v:5619" *) _T_4313;
  assign _T_4323 = _T_4297 ^ (* src = "crypto_accelerator.v:5620" *) _T_4295;
  assign _T_4325 = _T_4301 ^ (* src = "crypto_accelerator.v:5621" *) _T_4240;
  assign _T_4327 = _T_4307 ^ (* src = "crypto_accelerator.v:5622" *) _T_4305;
  assign _T_4329 = _T_4311 ^ (* src = "crypto_accelerator.v:5623" *) _T_4321;
  assign _T_4331 = _T_4323 ^ (* src = "crypto_accelerator.v:5624" *) _T_4317;
  assign _T_4333 = _T_4325 ^ (* src = "crypto_accelerator.v:5625" *) _T_4321;
  assign _T_4335 = _T_4327 ^ (* src = "crypto_accelerator.v:5626" *) _T_4317;
  assign _T_4337 = _T_4329 ^ (* src = "crypto_accelerator.v:5627" *) _T_4259;
  assign _T_4339 = _T_4335 ^ (* src = "crypto_accelerator.v:5628" *) _T_4337;
  assign _T_4343 = _T_4333 ^ (* src = "crypto_accelerator.v:5630" *) _T_4341;
  assign _T_4345 = _T_4331 ^ (* src = "crypto_accelerator.v:5631" *) _T_4333;
  assign _T_4347 = _T_4337 ^ (* src = "crypto_accelerator.v:5632" *) _T_4341;
  assign _T_4357 = _T_4345 ^ (* src = "crypto_accelerator.v:5637" *) _T_4341;
  assign _T_4363 = _T_4339 ^ (* src = "crypto_accelerator.v:5640" *) _T_4341;
  assign _T_4365 = _T_4333 ^ (* src = "crypto_accelerator.v:5641" *) _T_4349;
  assign _T_4367 = _T_4355 ^ (* src = "crypto_accelerator.v:5642" *) _T_4357;
  assign _T_4369 = _T_4337 ^ (* src = "crypto_accelerator.v:5643" *) _T_4351;
  assign _T_4371 = _T_4361 ^ (* src = "crypto_accelerator.v:5644" *) _T_4363;
  assign _T_4373 = _T_4367 ^ (* src = "crypto_accelerator.v:5645" *) _T_4371;
  assign _T_4375 = _T_4365 ^ (* src = "crypto_accelerator.v:5646" *) _T_4369;
  assign _T_4377 = _T_4365 ^ (* src = "crypto_accelerator.v:5647" *) _T_4367;
  assign _T_4379 = _T_4369 ^ (* src = "crypto_accelerator.v:5648" *) _T_4371;
  assign _T_4381 = _T_4375 ^ (* src = "crypto_accelerator.v:5649" *) _T_4373;
  assign _T_4419 = _T_4395 ^ (* src = "crypto_accelerator.v:5668" *) _T_4413;
  assign _T_4421 = _T_4407 ^ (* src = "crypto_accelerator.v:5669" *) _T_4409;
  assign _T_4423 = _T_4399 ^ (* src = "crypto_accelerator.v:5670" *) _T_4415;
  assign _T_4425 = _T_4385 ^ (* src = "crypto_accelerator.v:5671" *) _T_4391;
  assign _T_4427 = _T_4387 ^ (* src = "crypto_accelerator.v:5672" *) _T_4403;
  assign _T_4429 = _T_4383 ^ (* src = "crypto_accelerator.v:5673" *) _T_4393;
  assign _T_4431 = _T_4389 ^ (* src = "crypto_accelerator.v:5674" *) _T_4411;
  assign _T_4433 = _T_4419 ^ (* src = "crypto_accelerator.v:5675" *) _T_4421;
  assign _T_4435 = _T_4391 ^ (* src = "crypto_accelerator.v:5676" *) _T_4397;
  assign _T_4437 = _T_4401 ^ (* src = "crypto_accelerator.v:5677" *) _T_4417;
  assign _T_4439 = _T_4405 ^ (* src = "crypto_accelerator.v:5678" *) _T_4427;
  assign _T_4441 = _T_4419 ^ (* src = "crypto_accelerator.v:5679" *) _T_4425;
  assign _T_4443 = _T_4383 ^ (* src = "crypto_accelerator.v:5680" *) _T_4387;
  assign _T_4445 = _T_4389 ^ (* src = "crypto_accelerator.v:5681" *) _T_4393;
  assign _T_4447 = _T_4389 ^ (* src = "crypto_accelerator.v:5682" *) _T_4415;
  assign _T_4449 = _T_4399 ^ (* src = "crypto_accelerator.v:5683" *) _T_4409;
  assign _T_4451 = _T_4405 ^ (* src = "crypto_accelerator.v:5684" *) _T_4413;
  assign _T_4453 = _T_4407 ^ (* src = "crypto_accelerator.v:5685" *) _T_4423;
  assign _T_4455 = _T_4417 ^ (* src = "crypto_accelerator.v:5686" *) _T_4429;
  assign _T_4457 = _T_4423 ^ (* src = "crypto_accelerator.v:5687" *) _T_4425;
  assign _T_4459 = _T_4427 ^ (* src = "crypto_accelerator.v:5688" *) _T_4431;
  assign _T_4461 = _T_4423 ^ (* src = "crypto_accelerator.v:5689" *) _T_4433;
  assign _T_4463 = _T_4433 ^ (* src = "crypto_accelerator.v:5690" *) _T_4435;
  assign _T_4465 = _T_4429 ^ (* src = "crypto_accelerator.v:5691" *) _T_4433;
  assign _T_4467 = _T_4431 ^ (* src = "crypto_accelerator.v:5692" *) _T_4439;
  assign _T_4469 = _T_4437 ^ (* src = "crypto_accelerator.v:5693" *) _T_4441;
  assign _T_4471 = _T_4439 ^ (* src = "crypto_accelerator.v:5694" *) _T_4455;
  assign _T_4473 = _T_4441 ^ (* src = "crypto_accelerator.v:5695" *) _T_4467;
  assign _T_4475 = _T_4449 ^ (* src = "crypto_accelerator.v:5696" *) _T_4459;
  assign _T_4476 = _T_4445 ^ (* src = "crypto_accelerator.v:5697" *) _T_4461;
  assign _T_4477 = _T_4469 ^ (* src = "crypto_accelerator.v:5698" *) _T_4475;
  assign _T_4478 = _T_4453 ^ (* src = "crypto_accelerator.v:5699" *) _T_4473;
  assign _T_4479 = _T_4443 ^ (* src = "crypto_accelerator.v:5700" *) _T_4461;
  assign _T_4480 = _T_4463 ^ (* src = "crypto_accelerator.v:5701" *) _T_4471;
  assign _T_4481 = _T_4457 ^ (* src = "crypto_accelerator.v:5702" *) _T_4465;
  assign _T_4482 = _T_4447 ^ (* src = "crypto_accelerator.v:5703" *) _T_4463;
  assign _T_4483 = _T_4437 ^ (* src = "crypto_accelerator.v:5704" *) _T_4451;
  assign xorOut_0_0 = matrix_0_0 ^ (* src = "crypto_accelerator.v:5931" *) _GEN_224;
  assign xorOut_0_1 = matrix_0_1 ^ (* src = "crypto_accelerator.v:5932" *) _GEN_225;
  assign xorOut_0_2 = matrix_0_2 ^ (* src = "crypto_accelerator.v:5933" *) _GEN_226;
  assign xorOut_0_3 = matrix_0_3 ^ (* src = "crypto_accelerator.v:5934" *) _GEN_227;
  assign xorOut_1_0 = matrix_1_0 ^ (* src = "crypto_accelerator.v:5935" *) _GEN_228;
  assign xorOut_1_1 = matrix_1_1 ^ (* src = "crypto_accelerator.v:5936" *) _GEN_229;
  assign xorOut_1_2 = matrix_1_2 ^ (* src = "crypto_accelerator.v:5937" *) _GEN_230;
  assign xorOut_1_3 = matrix_1_3 ^ (* src = "crypto_accelerator.v:5938" *) _GEN_231;
  assign xorOut_2_0 = matrix_2_0 ^ (* src = "crypto_accelerator.v:5939" *) _GEN_232;
  assign xorOut_2_1 = matrix_2_1 ^ (* src = "crypto_accelerator.v:5940" *) _GEN_233;
  assign xorOut_2_2 = matrix_2_2 ^ (* src = "crypto_accelerator.v:5941" *) _GEN_234;
  assign xorOut_2_3 = matrix_2_3 ^ (* src = "crypto_accelerator.v:5942" *) _GEN_235;
  assign xorOut_3_0 = matrix_3_0 ^ (* src = "crypto_accelerator.v:5943" *) _GEN_236;
  assign xorOut_3_1 = matrix_3_1 ^ (* src = "crypto_accelerator.v:5944" *) _GEN_237;
  assign xorOut_3_2 = matrix_3_2 ^ (* src = "crypto_accelerator.v:5945" *) _GEN_238;
  assign xorOut_3_3 = matrix_3_3 ^ (* src = "crypto_accelerator.v:5946" *) _GEN_239;
  assign _T_4534 = xorOut_0_0 ^ (* src = "crypto_accelerator.v:5947" *) xorOut_0_2;
  assign _T_4538 = { _T_4534, 1'b0 } ^ (* src = "crypto_accelerator.v:5951" *) 5'b11011;
  assign _T_4545 = { _T_4541[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:5957" *) 5'b11011;
  assign _T_4549 = xorOut_0_1 ^ (* src = "crypto_accelerator.v:5960" *) xorOut_0_3;
  assign _T_4553 = { _T_4549, 1'b0 } ^ (* src = "crypto_accelerator.v:5964" *) 5'b11011;
  assign _T_4560 = { _T_4556[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:5970" *) 5'b11011;
  assign MixColsModule_io_in_0_0 = xorOut_0_0 ^ (* src = "crypto_accelerator.v:5974" *) _T_4548;
  assign MixColsModule_io_in_0_1 = xorOut_0_1 ^ (* src = "crypto_accelerator.v:5976" *) _T_4563;
  assign MixColsModule_io_in_0_2 = xorOut_0_2 ^ (* src = "crypto_accelerator.v:5978" *) _T_4548;
  assign MixColsModule_io_in_0_3 = xorOut_0_3 ^ (* src = "crypto_accelerator.v:5980" *) _T_4563;
  assign _T_4568 = xorOut_1_0 ^ (* src = "crypto_accelerator.v:5981" *) xorOut_1_2;
  assign _T_4572 = { _T_4568, 1'b0 } ^ (* src = "crypto_accelerator.v:5985" *) 5'b11011;
  assign _T_4579 = { _T_4575[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:5991" *) 5'b11011;
  assign _T_4583 = xorOut_1_1 ^ (* src = "crypto_accelerator.v:5994" *) xorOut_1_3;
  assign _T_4587 = { _T_4583, 1'b0 } ^ (* src = "crypto_accelerator.v:5998" *) 5'b11011;
  assign _T_4594 = { _T_4590[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:6004" *) 5'b11011;
  assign MixColsModule_io_in_1_0 = xorOut_1_0 ^ (* src = "crypto_accelerator.v:6008" *) _T_4582[7:0];
  assign MixColsModule_io_in_1_1 = xorOut_1_1 ^ (* src = "crypto_accelerator.v:6010" *) _T_4597;
  assign MixColsModule_io_in_1_2 = xorOut_1_2 ^ (* src = "crypto_accelerator.v:6012" *) _T_4582[7:0];
  assign MixColsModule_io_in_1_3 = xorOut_1_3 ^ (* src = "crypto_accelerator.v:6014" *) _T_4597;
  assign _T_4602 = xorOut_2_0 ^ (* src = "crypto_accelerator.v:6015" *) xorOut_2_2;
  assign _T_4606 = { _T_4602, 1'b0 } ^ (* src = "crypto_accelerator.v:6019" *) 5'b11011;
  assign _T_4613 = { _T_4609[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:6025" *) 5'b11011;
  assign _T_4617 = xorOut_2_1 ^ (* src = "crypto_accelerator.v:6028" *) xorOut_2_3;
  assign _T_4621 = { _T_4617, 1'b0 } ^ (* src = "crypto_accelerator.v:6032" *) 5'b11011;
  assign _T_4628 = { _T_4624[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:6038" *) 5'b11011;
  assign MixColsModule_io_in_2_0 = xorOut_2_0 ^ (* src = "crypto_accelerator.v:6042" *) _T_4616[7:0];
  assign MixColsModule_io_in_2_1 = xorOut_2_1 ^ (* src = "crypto_accelerator.v:6044" *) _T_4631[7:0];
  assign MixColsModule_io_in_2_2 = xorOut_2_2 ^ (* src = "crypto_accelerator.v:6046" *) _T_4616[7:0];
  assign MixColsModule_io_in_2_3 = xorOut_2_3 ^ (* src = "crypto_accelerator.v:6048" *) _T_4631[7:0];
  assign _T_4636 = xorOut_3_0 ^ (* src = "crypto_accelerator.v:6049" *) xorOut_3_2;
  assign _T_4640 = { _T_4636, 1'b0 } ^ (* src = "crypto_accelerator.v:6053" *) 5'b11011;
  assign _T_4647 = { _T_4643[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:6059" *) 5'b11011;
  assign _T_4651 = xorOut_3_1 ^ (* src = "crypto_accelerator.v:6062" *) xorOut_3_3;
  assign _T_4655 = { _T_4651, 1'b0 } ^ (* src = "crypto_accelerator.v:6066" *) 5'b11011;
  assign _T_4662 = { _T_4658[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:6072" *) 5'b11011;
  assign MixColsModule_io_in_3_0 = xorOut_3_0 ^ (* src = "crypto_accelerator.v:6076" *) _T_4650[7:0];
  assign MixColsModule_io_in_3_1 = xorOut_3_1 ^ (* src = "crypto_accelerator.v:6078" *) _T_4665;
  assign MixColsModule_io_in_3_2 = xorOut_3_2 ^ (* src = "crypto_accelerator.v:6080" *) _T_4650[7:0];
  assign MixColsModule_io_in_3_3 = xorOut_3_3 ^ (* src = "crypto_accelerator.v:6082" *) _T_4665;
  assign _T_4726 = io_ivIn ^ (* src = "crypto_accelerator.v:6085" *) { xorOut_0_0, xorOut_0_1, xorOut_0_2, xorOut_0_3, xorOut_1_0, xorOut_1_1, xorOut_1_2, xorOut_1_3, xorOut_2_0, xorOut_2_1, xorOut_2_2, xorOut_2_3, xorOut_3_0, xorOut_3_1, xorOut_3_2, xorOut_3_3 };
  (* src = "crypto_accelerator.v:6112" *)
  MixColsModule MixColsModule (
    .io_in_0_0(MixColsModule_io_in_0_0),
    .io_in_0_1(MixColsModule_io_in_0_1),
    .io_in_0_2(MixColsModule_io_in_0_2),
    .io_in_0_3(MixColsModule_io_in_0_3),
    .io_in_1_0(MixColsModule_io_in_1_0),
    .io_in_1_1(MixColsModule_io_in_1_1),
    .io_in_1_2(MixColsModule_io_in_1_2),
    .io_in_1_3(MixColsModule_io_in_1_3),
    .io_in_2_0(MixColsModule_io_in_2_0),
    .io_in_2_1(MixColsModule_io_in_2_1),
    .io_in_2_2(MixColsModule_io_in_2_2),
    .io_in_2_3(MixColsModule_io_in_2_3),
    .io_in_3_0(MixColsModule_io_in_3_0),
    .io_in_3_1(MixColsModule_io_in_3_1),
    .io_in_3_2(MixColsModule_io_in_3_2),
    .io_in_3_3(MixColsModule_io_in_3_3),
    .io_out_0_0(MixColsModule_io_out_0_0),
    .io_out_0_1(MixColsModule_io_out_0_1),
    .io_out_0_2(MixColsModule_io_out_0_2),
    .io_out_0_3(MixColsModule_io_out_0_3),
    .io_out_1_0(MixColsModule_io_out_1_0),
    .io_out_1_1(MixColsModule_io_out_1_1),
    .io_out_1_2(MixColsModule_io_out_1_2),
    .io_out_1_3(MixColsModule_io_out_1_3),
    .io_out_2_0(MixColsModule_io_out_2_0),
    .io_out_2_1(MixColsModule_io_out_2_1),
    .io_out_2_2(MixColsModule_io_out_2_2),
    .io_out_2_3(MixColsModule_io_out_2_3),
    .io_out_3_0(MixColsModule_io_out_3_0),
    .io_out_3_1(MixColsModule_io_out_3_1),
    .io_out_3_2(MixColsModule_io_out_3_2),
    .io_out_3_3(MixColsModule_io_out_3_3)
  );
  assign _GEN_100 = io_keys_0_1_0;
  assign _GEN_101 = io_keys_0_1_1;
  assign _GEN_102 = io_keys_0_1_2;
  assign _GEN_103 = io_keys_0_1_3;
  assign _GEN_104 = io_keys_0_2_0;
  assign _GEN_105 = io_keys_0_2_1;
  assign _GEN_106 = io_keys_0_2_2;
  assign _GEN_107 = io_keys_0_2_3;
  assign _GEN_108 = io_keys_0_3_0;
  assign _GEN_109 = io_keys_0_3_1;
  assign _GEN_110 = io_keys_0_3_2;
  assign _GEN_111 = io_keys_0_3_3;
  assign _GEN_112 = io_keys_0_0_0;
  assign _GEN_113 = io_keys_0_0_1;
  assign _GEN_114 = io_keys_0_0_2;
  assign _GEN_115 = io_keys_0_0_3;
  assign _GEN_116 = io_keys_0_1_0;
  assign _GEN_117 = io_keys_0_1_1;
  assign _GEN_118 = io_keys_0_1_2;
  assign _GEN_119 = io_keys_0_1_3;
  assign _GEN_120 = io_keys_0_2_0;
  assign _GEN_121 = io_keys_0_2_1;
  assign _GEN_122 = io_keys_0_2_2;
  assign _GEN_123 = io_keys_0_2_3;
  assign _GEN_124 = io_keys_0_3_0;
  assign _GEN_125 = io_keys_0_3_1;
  assign _GEN_126 = io_keys_0_3_2;
  assign _GEN_127 = io_keys_0_3_3;
  assign _GEN_16 = io_keys_0_0_0;
  assign _GEN_17 = io_keys_0_0_1;
  assign _GEN_18 = io_keys_0_0_2;
  assign _GEN_19 = io_keys_0_0_3;
  assign _GEN_20 = io_keys_0_1_0;
  assign _GEN_21 = io_keys_0_1_1;
  assign _GEN_22 = io_keys_0_1_2;
  assign _GEN_23 = io_keys_0_1_3;
  assign _GEN_24 = io_keys_0_2_0;
  assign _GEN_25 = io_keys_0_2_1;
  assign _GEN_26 = io_keys_0_2_2;
  assign _GEN_27 = io_keys_0_2_3;
  assign _GEN_275 = state[0];
  assign _GEN_28 = io_keys_0_3_0;
  assign _GEN_29 = io_keys_0_3_1;
  assign _GEN_30 = io_keys_0_3_2;
  assign _GEN_31 = io_keys_0_3_3;
  assign _GEN_311 = { 2'b00, xorOut_0_0 };
  assign _GEN_312 = { 2'b00, xorOut_0_1 };
  assign _GEN_313 = { 2'b00, xorOut_0_2 };
  assign _GEN_314 = { 2'b00, xorOut_0_3 };
  assign _GEN_315 = { 2'b00, xorOut_1_0 };
  assign _GEN_316 = { 2'b00, xorOut_1_1 };
  assign _GEN_317 = { 2'b00, xorOut_1_2 };
  assign _GEN_318 = { 2'b00, xorOut_1_3 };
  assign _GEN_319 = { 2'b00, xorOut_2_0 };
  assign _GEN_32 = io_keys_0_0_0;
  assign _GEN_320 = { 2'b00, xorOut_2_1 };
  assign _GEN_321 = { 2'b00, xorOut_2_2 };
  assign _GEN_322 = { 2'b00, xorOut_2_3 };
  assign _GEN_323 = { 2'b00, xorOut_3_0 };
  assign _GEN_324 = { 2'b00, xorOut_3_1 };
  assign _GEN_325 = { 2'b00, xorOut_3_2 };
  assign _GEN_326 = { 2'b00, xorOut_3_3 };
  assign _GEN_33 = io_keys_0_0_1;
  assign _GEN_34 = io_keys_0_0_2;
  assign _GEN_35 = io_keys_0_0_3;
  assign _GEN_36 = io_keys_0_1_0;
  assign _GEN_37 = io_keys_0_1_1;
  assign _GEN_38 = io_keys_0_1_2;
  assign _GEN_39 = io_keys_0_1_3;
  assign _GEN_40 = io_keys_0_2_0;
  assign _GEN_41 = io_keys_0_2_1;
  assign _GEN_42 = io_keys_0_2_2;
  assign _GEN_43 = io_keys_0_2_3;
  assign _GEN_44 = io_keys_0_3_0;
  assign _GEN_45 = io_keys_0_3_1;
  assign _GEN_46 = io_keys_0_3_2;
  assign _GEN_47 = io_keys_0_3_3;
  assign _GEN_48 = io_keys_0_0_0;
  assign _GEN_49 = io_keys_0_0_1;
  assign _GEN_50 = io_keys_0_0_2;
  assign _GEN_51 = io_keys_0_0_3;
  assign _GEN_52 = io_keys_0_1_0;
  assign _GEN_53 = io_keys_0_1_1;
  assign _GEN_54 = io_keys_0_1_2;
  assign _GEN_55 = io_keys_0_1_3;
  assign _GEN_56 = io_keys_0_2_0;
  assign _GEN_57 = io_keys_0_2_1;
  assign _GEN_58 = io_keys_0_2_2;
  assign _GEN_59 = io_keys_0_2_3;
  assign _GEN_60 = io_keys_0_3_0;
  assign _GEN_61 = io_keys_0_3_1;
  assign _GEN_62 = io_keys_0_3_2;
  assign _GEN_63 = io_keys_0_3_3;
  assign _GEN_64 = io_keys_0_0_0;
  assign _GEN_65 = io_keys_0_0_1;
  assign _GEN_66 = io_keys_0_0_2;
  assign _GEN_67 = io_keys_0_0_3;
  assign _GEN_68 = io_keys_0_1_0;
  assign _GEN_69 = io_keys_0_1_1;
  assign _GEN_70 = io_keys_0_1_2;
  assign _GEN_71 = io_keys_0_1_3;
  assign _GEN_72 = io_keys_0_2_0;
  assign _GEN_73 = io_keys_0_2_1;
  assign _GEN_74 = io_keys_0_2_2;
  assign _GEN_75 = io_keys_0_2_3;
  assign _GEN_76 = io_keys_0_3_0;
  assign _GEN_77 = io_keys_0_3_1;
  assign _GEN_78 = io_keys_0_3_2;
  assign _GEN_79 = io_keys_0_3_3;
  assign _GEN_80 = io_keys_0_0_0;
  assign _GEN_81 = io_keys_0_0_1;
  assign _GEN_82 = io_keys_0_0_2;
  assign _GEN_83 = io_keys_0_0_3;
  assign _GEN_84 = io_keys_0_1_0;
  assign _GEN_85 = io_keys_0_1_1;
  assign _GEN_86 = io_keys_0_1_2;
  assign _GEN_87 = io_keys_0_1_3;
  assign _GEN_88 = io_keys_0_2_0;
  assign _GEN_89 = io_keys_0_2_1;
  assign _GEN_90 = io_keys_0_2_2;
  assign _GEN_91 = io_keys_0_2_3;
  assign _GEN_92 = io_keys_0_3_0;
  assign _GEN_93 = io_keys_0_3_1;
  assign _GEN_94 = io_keys_0_3_2;
  assign _GEN_95 = io_keys_0_3_3;
  assign _GEN_96 = io_keys_0_0_0;
  assign _GEN_97 = io_keys_0_0_1;
  assign _GEN_98 = io_keys_0_0_2;
  assign _GEN_99 = io_keys_0_0_3;
  assign _T_10 = { matrix_2_0, matrix_2_1, matrix_2_2, matrix_2_3, matrix_3_0, matrix_3_1, matrix_3_2, matrix_3_3 };
  assign _T_17 = { matrix_0_0, matrix_0_1, matrix_0_2, matrix_0_3, matrix_1_0, matrix_1_1, matrix_1_2, matrix_1_3 };
  assign _T_4537 = { _T_4534, 1'b0 };
  assign _T_4544 = { _T_4541, 1'b0 };
  assign _T_4552 = { _T_4549, 1'b0 };
  assign _T_4559 = { _T_4556, 1'b0 };
  assign _T_4564[7:0] = MixColsModule_io_in_0_0;
  assign _T_4565[7:0] = MixColsModule_io_in_0_1;
  assign _T_4566[7:0] = MixColsModule_io_in_0_2;
  assign _T_4567[7:0] = MixColsModule_io_in_0_3;
  assign _T_4571 = { _T_4568, 1'b0 };
  assign _T_4578 = { _T_4575, 1'b0 };
  assign _T_4582[9:8] = 2'bxx;
  assign _T_4586 = { _T_4583, 1'b0 };
  assign _T_4593 = { _T_4590, 1'b0 };
  assign _T_4598[7:0] = MixColsModule_io_in_1_0;
  assign _T_4599[7:0] = MixColsModule_io_in_1_1;
  assign _T_4600[7:0] = MixColsModule_io_in_1_2;
  assign _T_4601[7:0] = MixColsModule_io_in_1_3;
  assign _T_4605 = { _T_4602, 1'b0 };
  assign _T_4612 = { _T_4609, 1'b0 };
  assign _T_4616[9:8] = 2'bxx;
  assign _T_4620 = { _T_4617, 1'b0 };
  assign _T_4627 = { _T_4624, 1'b0 };
  assign _T_4631[9:8] = 2'bxx;
  assign _T_4632[7:0] = MixColsModule_io_in_2_0;
  assign _T_4633[7:0] = MixColsModule_io_in_2_1;
  assign _T_4634[7:0] = MixColsModule_io_in_2_2;
  assign _T_4635[7:0] = MixColsModule_io_in_2_3;
  assign _T_4639 = { _T_4636, 1'b0 };
  assign _T_4646 = { _T_4643, 1'b0 };
  assign _T_4650[9:8] = 2'bxx;
  assign _T_4654 = { _T_4651, 1'b0 };
  assign _T_4661 = { _T_4658, 1'b0 };
  assign _T_4666[7:0] = MixColsModule_io_in_3_0;
  assign _T_4667[7:0] = MixColsModule_io_in_3_1;
  assign _T_4668[7:0] = MixColsModule_io_in_3_2;
  assign _T_4669[7:0] = MixColsModule_io_in_3_3;
  assign _T_4717 = { xorOut_2_0, xorOut_2_1, xorOut_2_2, xorOut_2_3, xorOut_3_0, xorOut_3_1, xorOut_3_2, xorOut_3_3 };
  assign _T_4725 = { xorOut_0_0, xorOut_0_1, xorOut_0_2, xorOut_0_3, xorOut_1_0, xorOut_1_1, xorOut_1_2, xorOut_1_3, xorOut_2_0, xorOut_2_1, xorOut_2_2, xorOut_2_3, xorOut_3_0, xorOut_3_1, xorOut_3_2, xorOut_3_3 };
  assign _T_4769 = _GEN_327;
  assign finalOut_0_0 = _T_4726[127:120];
  assign finalOut_0_1 = _T_4726[119:112];
  assign finalOut_0_2 = _T_4726[111:104];
  assign finalOut_0_3 = _T_4726[103:96];
  assign finalOut_1_0 = _T_4726[95:88];
  assign finalOut_1_1 = _T_4726[87:80];
  assign finalOut_1_2 = _T_4726[79:72];
  assign finalOut_1_3 = _T_4726[71:64];
  assign finalOut_2_0 = _T_4726[63:56];
  assign finalOut_2_1 = _T_4726[55:48];
  assign finalOut_2_2 = _T_4726[47:40];
  assign finalOut_2_3 = _T_4726[39:32];
  assign finalOut_3_0 = _T_4726[31:24];
  assign finalOut_3_1 = _T_4726[23:16];
  assign finalOut_3_2 = _T_4726[15:8];
  assign finalOut_3_3 = _T_4726[7:0];
  assign io_dataOut = { matrix_0_0, matrix_0_1, matrix_0_2, matrix_0_3, matrix_1_0, matrix_1_1, matrix_1_2, matrix_1_3, matrix_2_0, matrix_2_1, matrix_2_2, matrix_2_3, matrix_3_0, matrix_3_1, matrix_3_2, matrix_3_3 };
  assign io_ivOut = ctSaved;
  assign io_outputValid = _T;
  assign io_shiftCyc = io_shift;
  assign io_shiftRev = io_shift;
  assign roundPart1_0_0 = { _T_288, _T_289, _T_290, _T_291, _T_292, _T_293, _T_294, _T_295 };
  assign roundPart1_0_1 = { _T_567, _T_568, _T_569, _T_570, _T_571, _T_572, _T_573, _T_574 };
  assign roundPart1_0_2 = { _T_846, _T_847, _T_848, _T_849, _T_850, _T_851, _T_852, _T_853 };
  assign roundPart1_0_3 = { _T_1125, _T_1126, _T_1127, _T_1128, _T_1129, _T_1130, _T_1131, _T_1132 };
  assign roundPart1_1_0 = { _T_1405, _T_1406, _T_1407, _T_1408, _T_1409, _T_1410, _T_1411, _T_1412 };
  assign roundPart1_1_1 = { _T_1684, _T_1685, _T_1686, _T_1687, _T_1688, _T_1689, _T_1690, _T_1691 };
  assign roundPart1_1_2 = { _T_1963, _T_1964, _T_1965, _T_1966, _T_1967, _T_1968, _T_1969, _T_1970 };
  assign roundPart1_1_3 = { _T_2242, _T_2243, _T_2244, _T_2245, _T_2246, _T_2247, _T_2248, _T_2249 };
  assign roundPart1_2_0 = { _T_2522, _T_2523, _T_2524, _T_2525, _T_2526, _T_2527, _T_2528, _T_2529 };
  assign roundPart1_2_1 = { _T_2801, _T_2802, _T_2803, _T_2804, _T_2805, _T_2806, _T_2807, _T_2808 };
  assign roundPart1_2_2 = { _T_3080, _T_3081, _T_3082, _T_3083, _T_3084, _T_3085, _T_3086, _T_3087 };
  assign roundPart1_2_3 = { _T_3359, _T_3360, _T_3361, _T_3362, _T_3363, _T_3364, _T_3365, _T_3366 };
  assign roundPart1_3_0 = { _T_3639, _T_3640, _T_3641, _T_3642, _T_3643, _T_3644, _T_3645, _T_3646 };
  assign roundPart1_3_1 = { _T_3918, _T_3919, _T_3920, _T_3921, _T_3922, _T_3923, _T_3924, _T_3925 };
  assign roundPart1_3_2 = { _T_4197, _T_4198, _T_4199, _T_4200, _T_4201, _T_4202, _T_4203, _T_4204 };
  assign roundPart1_3_3 = { _T_4476, _T_4477, _T_4478, _T_4479, _T_4480, _T_4481, _T_4482, _T_4483 };
endmodule
