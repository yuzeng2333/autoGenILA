module \$paramod\SDP_C_mgc_in_wire_v1\rscid=4\width=6 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:78" *)
  output [5:0] d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:79" *)
  input [5:0] z;
  assign d = z;
endmodule
