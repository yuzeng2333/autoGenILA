module ShiftRegister_1(clock, io_input, io_enable, io_output_1, io_output_6, io_output_14, io_output_15);
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _00_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _01_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _02_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _03_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _04_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _05_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _06_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _07_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _08_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _09_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _10_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _11_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _12_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _13_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _14_;
  (* src = "crypto_accelerator.v:8591" *)
  wire [31:0] _15_;
  (* src = "crypto_accelerator.v:8471" *)
  input clock;
  (* src = "crypto_accelerator.v:8473" *)
  input io_enable;
  (* src = "crypto_accelerator.v:8472" *)
  input [31:0] io_input;
  (* src = "crypto_accelerator.v:8474" *)
  output [31:0] io_output_1;
  (* src = "crypto_accelerator.v:8476" *)
  output [31:0] io_output_14;
  (* src = "crypto_accelerator.v:8477" *)
  output [31:0] io_output_15;
  (* src = "crypto_accelerator.v:8475" *)
  output [31:0] io_output_6;
  (* src = "crypto_accelerator.v:8497" *)
  reg [31:0] reg_0;
  (* src = "crypto_accelerator.v:8498" *)
  reg [31:0] reg_1;
  (* src = "crypto_accelerator.v:8507" *)
  reg [31:0] reg_10;
  (* src = "crypto_accelerator.v:8508" *)
  reg [31:0] reg_11;
  (* src = "crypto_accelerator.v:8509" *)
  reg [31:0] reg_12;
  (* src = "crypto_accelerator.v:8510" *)
  reg [31:0] reg_13;
  (* src = "crypto_accelerator.v:8511" *)
  reg [31:0] reg_14;
  (* src = "crypto_accelerator.v:8512" *)
  reg [31:0] reg_15;
  (* src = "crypto_accelerator.v:8499" *)
  reg [31:0] reg_2;
  (* src = "crypto_accelerator.v:8500" *)
  reg [31:0] reg_3;
  (* src = "crypto_accelerator.v:8501" *)
  reg [31:0] reg_4;
  (* src = "crypto_accelerator.v:8502" *)
  reg [31:0] reg_5;
  (* src = "crypto_accelerator.v:8503" *)
  reg [31:0] reg_6;
  (* src = "crypto_accelerator.v:8504" *)
  reg [31:0] reg_7;
  (* src = "crypto_accelerator.v:8505" *)
  reg [31:0] reg_8;
  (* src = "crypto_accelerator.v:8506" *)
  reg [31:0] reg_9;
  always @(posedge clock)
      reg_0 <= _00_;
  always @(posedge clock)
      reg_1 <= _07_;
  always @(posedge clock)
      reg_2 <= _08_;
  always @(posedge clock)
      reg_3 <= _09_;
  always @(posedge clock)
      reg_4 <= _10_;
  always @(posedge clock)
      reg_5 <= _11_;
  always @(posedge clock)
      reg_6 <= _12_;
  always @(posedge clock)
      reg_7 <= _13_;
  always @(posedge clock)
      reg_8 <= _14_;
  always @(posedge clock)
      reg_9 <= _15_;
  always @(posedge clock)
      reg_10 <= _01_;
  always @(posedge clock)
      reg_11 <= _02_;
  always @(posedge clock)
      reg_12 <= _03_;
  always @(posedge clock)
      reg_13 <= _04_;
  always @(posedge clock)
      reg_14 <= _05_;
  always @(posedge clock)
      reg_15 <= _06_;
  assign _06_ = io_enable ? (* src = "crypto_accelerator.v:8637" *) reg_14 : reg_15;
  assign _05_ = io_enable ? (* src = "crypto_accelerator.v:8634" *) reg_13 : reg_14;
  assign _04_ = io_enable ? (* src = "crypto_accelerator.v:8631" *) reg_12 : reg_13;
  assign _03_ = io_enable ? (* src = "crypto_accelerator.v:8628" *) reg_11 : reg_12;
  assign _02_ = io_enable ? (* src = "crypto_accelerator.v:8625" *) reg_10 : reg_11;
  assign _01_ = io_enable ? (* src = "crypto_accelerator.v:8622" *) reg_9 : reg_10;
  assign _15_ = io_enable ? (* src = "crypto_accelerator.v:8619" *) reg_8 : reg_9;
  assign _14_ = io_enable ? (* src = "crypto_accelerator.v:8616" *) reg_7 : reg_8;
  assign _13_ = io_enable ? (* src = "crypto_accelerator.v:8613" *) reg_6 : reg_7;
  assign _12_ = io_enable ? (* src = "crypto_accelerator.v:8610" *) reg_5 : reg_6;
  assign _11_ = io_enable ? (* src = "crypto_accelerator.v:8607" *) reg_4 : reg_5;
  assign _10_ = io_enable ? (* src = "crypto_accelerator.v:8604" *) reg_3 : reg_4;
  assign _09_ = io_enable ? (* src = "crypto_accelerator.v:8601" *) reg_2 : reg_3;
  assign _08_ = io_enable ? (* src = "crypto_accelerator.v:8598" *) reg_1 : reg_2;
  assign _07_ = io_enable ? (* src = "crypto_accelerator.v:8595" *) reg_0 : reg_1;
  assign _00_ = io_enable ? (* src = "crypto_accelerator.v:8592" *) io_input : reg_0;
  assign io_output_1 = reg_1;
  assign io_output_14 = reg_14;
  assign io_output_15 = reg_15;
  assign io_output_6 = reg_6;
endmodule
