module \$paramod\CSC_mgc_in_wire_v1\rscid=3\width=2 (d, z);
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:78" *)
  output [1:0] d;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:79" *)
  input [1:0] z;
  assign d = z;
endmodule
