module NV_NVDLA_RT_csc2cmac_b(nvdla_core_clk, nvdla_core_rstn, sc2mac_wt_src_pvld, sc2mac_wt_src_mask, sc2mac_wt_src_data0, sc2mac_wt_src_data1, sc2mac_wt_src_data2, sc2mac_wt_src_data3, sc2mac_wt_src_data4, sc2mac_wt_src_data5, sc2mac_wt_src_data6, sc2mac_wt_src_data7, sc2mac_wt_src_data8, sc2mac_wt_src_data9, sc2mac_wt_src_data10, sc2mac_wt_src_data11, sc2mac_wt_src_data12, sc2mac_wt_src_data13, sc2mac_wt_src_data14, sc2mac_wt_src_data15, sc2mac_wt_src_data16, sc2mac_wt_src_data17, sc2mac_wt_src_data18, sc2mac_wt_src_data19, sc2mac_wt_src_data20, sc2mac_wt_src_data21, sc2mac_wt_src_data22, sc2mac_wt_src_data23, sc2mac_wt_src_data24, sc2mac_wt_src_data25, sc2mac_wt_src_data26, sc2mac_wt_src_data27, sc2mac_wt_src_data28, sc2mac_wt_src_data29, sc2mac_wt_src_data30, sc2mac_wt_src_data31, sc2mac_wt_src_data32, sc2mac_wt_src_data33, sc2mac_wt_src_data34, sc2mac_wt_src_data35, sc2mac_wt_src_data36, sc2mac_wt_src_data37, sc2mac_wt_src_data38, sc2mac_wt_src_data39, sc2mac_wt_src_data40, sc2mac_wt_src_data41, sc2mac_wt_src_data42, sc2mac_wt_src_data43, sc2mac_wt_src_data44, sc2mac_wt_src_data45, sc2mac_wt_src_data46, sc2mac_wt_src_data47, sc2mac_wt_src_data48, sc2mac_wt_src_data49, sc2mac_wt_src_data50, sc2mac_wt_src_data51, sc2mac_wt_src_data52, sc2mac_wt_src_data53, sc2mac_wt_src_data54, sc2mac_wt_src_data55, sc2mac_wt_src_data56, sc2mac_wt_src_data57, sc2mac_wt_src_data58, sc2mac_wt_src_data59, sc2mac_wt_src_data60, sc2mac_wt_src_data61, sc2mac_wt_src_data62, sc2mac_wt_src_data63, sc2mac_wt_src_data64, sc2mac_wt_src_data65, sc2mac_wt_src_data66, sc2mac_wt_src_data67, sc2mac_wt_src_data68, sc2mac_wt_src_data69, sc2mac_wt_src_data70, sc2mac_wt_src_data71, sc2mac_wt_src_data72, sc2mac_wt_src_data73, sc2mac_wt_src_data74, sc2mac_wt_src_data75, sc2mac_wt_src_data76, sc2mac_wt_src_data77, sc2mac_wt_src_data78, sc2mac_wt_src_data79, sc2mac_wt_src_data80, sc2mac_wt_src_data81, sc2mac_wt_src_data82, sc2mac_wt_src_data83, sc2mac_wt_src_data84, sc2mac_wt_src_data85, sc2mac_wt_src_data86, sc2mac_wt_src_data87, sc2mac_wt_src_data88, sc2mac_wt_src_data89, sc2mac_wt_src_data90, sc2mac_wt_src_data91, sc2mac_wt_src_data92, sc2mac_wt_src_data93, sc2mac_wt_src_data94, sc2mac_wt_src_data95, sc2mac_wt_src_data96, sc2mac_wt_src_data97, sc2mac_wt_src_data98, sc2mac_wt_src_data99, sc2mac_wt_src_data100, sc2mac_wt_src_data101, sc2mac_wt_src_data102, sc2mac_wt_src_data103, sc2mac_wt_src_data104, sc2mac_wt_src_data105, sc2mac_wt_src_data106, sc2mac_wt_src_data107, sc2mac_wt_src_data108, sc2mac_wt_src_data109, sc2mac_wt_src_data110, sc2mac_wt_src_data111, sc2mac_wt_src_data112, sc2mac_wt_src_data113, sc2mac_wt_src_data114, sc2mac_wt_src_data115, sc2mac_wt_src_data116, sc2mac_wt_src_data117, sc2mac_wt_src_data118, sc2mac_wt_src_data119, sc2mac_wt_src_data120, sc2mac_wt_src_data121, sc2mac_wt_src_data122, sc2mac_wt_src_data123, sc2mac_wt_src_data124, sc2mac_wt_src_data125, sc2mac_wt_src_data126, sc2mac_wt_src_data127, sc2mac_wt_src_sel, sc2mac_dat_src_pvld, sc2mac_dat_src_mask, sc2mac_dat_src_data0, sc2mac_dat_src_data1, sc2mac_dat_src_data2, sc2mac_dat_src_data3, sc2mac_dat_src_data4, sc2mac_dat_src_data5, sc2mac_dat_src_data6, sc2mac_dat_src_data7, sc2mac_dat_src_data8, sc2mac_dat_src_data9, sc2mac_dat_src_data10, sc2mac_dat_src_data11, sc2mac_dat_src_data12, sc2mac_dat_src_data13, sc2mac_dat_src_data14, sc2mac_dat_src_data15, sc2mac_dat_src_data16, sc2mac_dat_src_data17, sc2mac_dat_src_data18, sc2mac_dat_src_data19, sc2mac_dat_src_data20, sc2mac_dat_src_data21, sc2mac_dat_src_data22, sc2mac_dat_src_data23, sc2mac_dat_src_data24, sc2mac_dat_src_data25, sc2mac_dat_src_data26, sc2mac_dat_src_data27, sc2mac_dat_src_data28, sc2mac_dat_src_data29, sc2mac_dat_src_data30, sc2mac_dat_src_data31, sc2mac_dat_src_data32, sc2mac_dat_src_data33, sc2mac_dat_src_data34, sc2mac_dat_src_data35, sc2mac_dat_src_data36, sc2mac_dat_src_data37, sc2mac_dat_src_data38, sc2mac_dat_src_data39, sc2mac_dat_src_data40, sc2mac_dat_src_data41, sc2mac_dat_src_data42, sc2mac_dat_src_data43, sc2mac_dat_src_data44, sc2mac_dat_src_data45, sc2mac_dat_src_data46, sc2mac_dat_src_data47, sc2mac_dat_src_data48, sc2mac_dat_src_data49, sc2mac_dat_src_data50, sc2mac_dat_src_data51, sc2mac_dat_src_data52, sc2mac_dat_src_data53, sc2mac_dat_src_data54, sc2mac_dat_src_data55, sc2mac_dat_src_data56, sc2mac_dat_src_data57, sc2mac_dat_src_data58, sc2mac_dat_src_data59, sc2mac_dat_src_data60, sc2mac_dat_src_data61, sc2mac_dat_src_data62, sc2mac_dat_src_data63, sc2mac_dat_src_data64, sc2mac_dat_src_data65, sc2mac_dat_src_data66, sc2mac_dat_src_data67, sc2mac_dat_src_data68, sc2mac_dat_src_data69, sc2mac_dat_src_data70, sc2mac_dat_src_data71, sc2mac_dat_src_data72, sc2mac_dat_src_data73, sc2mac_dat_src_data74, sc2mac_dat_src_data75, sc2mac_dat_src_data76, sc2mac_dat_src_data77, sc2mac_dat_src_data78, sc2mac_dat_src_data79, sc2mac_dat_src_data80, sc2mac_dat_src_data81, sc2mac_dat_src_data82, sc2mac_dat_src_data83, sc2mac_dat_src_data84, sc2mac_dat_src_data85, sc2mac_dat_src_data86, sc2mac_dat_src_data87, sc2mac_dat_src_data88, sc2mac_dat_src_data89, sc2mac_dat_src_data90, sc2mac_dat_src_data91, sc2mac_dat_src_data92, sc2mac_dat_src_data93, sc2mac_dat_src_data94, sc2mac_dat_src_data95, sc2mac_dat_src_data96, sc2mac_dat_src_data97, sc2mac_dat_src_data98, sc2mac_dat_src_data99, sc2mac_dat_src_data100, sc2mac_dat_src_data101, sc2mac_dat_src_data102, sc2mac_dat_src_data103, sc2mac_dat_src_data104, sc2mac_dat_src_data105, sc2mac_dat_src_data106, sc2mac_dat_src_data107, sc2mac_dat_src_data108, sc2mac_dat_src_data109, sc2mac_dat_src_data110, sc2mac_dat_src_data111, sc2mac_dat_src_data112, sc2mac_dat_src_data113, sc2mac_dat_src_data114, sc2mac_dat_src_data115, sc2mac_dat_src_data116, sc2mac_dat_src_data117, sc2mac_dat_src_data118, sc2mac_dat_src_data119, sc2mac_dat_src_data120, sc2mac_dat_src_data121, sc2mac_dat_src_data122, sc2mac_dat_src_data123, sc2mac_dat_src_data124, sc2mac_dat_src_data125, sc2mac_dat_src_data126, sc2mac_dat_src_data127, sc2mac_dat_src_pd, sc2mac_wt_dst_pvld, sc2mac_wt_dst_mask, sc2mac_wt_dst_data0, sc2mac_wt_dst_data1, sc2mac_wt_dst_data2, sc2mac_wt_dst_data3, sc2mac_wt_dst_data4, sc2mac_wt_dst_data5, sc2mac_wt_dst_data6, sc2mac_wt_dst_data7, sc2mac_wt_dst_data8, sc2mac_wt_dst_data9, sc2mac_wt_dst_data10, sc2mac_wt_dst_data11, sc2mac_wt_dst_data12, sc2mac_wt_dst_data13, sc2mac_wt_dst_data14, sc2mac_wt_dst_data15, sc2mac_wt_dst_data16, sc2mac_wt_dst_data17, sc2mac_wt_dst_data18, sc2mac_wt_dst_data19, sc2mac_wt_dst_data20, sc2mac_wt_dst_data21, sc2mac_wt_dst_data22, sc2mac_wt_dst_data23, sc2mac_wt_dst_data24, sc2mac_wt_dst_data25, sc2mac_wt_dst_data26, sc2mac_wt_dst_data27, sc2mac_wt_dst_data28, sc2mac_wt_dst_data29, sc2mac_wt_dst_data30, sc2mac_wt_dst_data31, sc2mac_wt_dst_data32, sc2mac_wt_dst_data33, sc2mac_wt_dst_data34, sc2mac_wt_dst_data35, sc2mac_wt_dst_data36, sc2mac_wt_dst_data37, sc2mac_wt_dst_data38, sc2mac_wt_dst_data39, sc2mac_wt_dst_data40, sc2mac_wt_dst_data41, sc2mac_wt_dst_data42, sc2mac_wt_dst_data43, sc2mac_wt_dst_data44, sc2mac_wt_dst_data45, sc2mac_wt_dst_data46, sc2mac_wt_dst_data47, sc2mac_wt_dst_data48, sc2mac_wt_dst_data49, sc2mac_wt_dst_data50, sc2mac_wt_dst_data51, sc2mac_wt_dst_data52, sc2mac_wt_dst_data53, sc2mac_wt_dst_data54, sc2mac_wt_dst_data55, sc2mac_wt_dst_data56, sc2mac_wt_dst_data57, sc2mac_wt_dst_data58, sc2mac_wt_dst_data59, sc2mac_wt_dst_data60, sc2mac_wt_dst_data61, sc2mac_wt_dst_data62, sc2mac_wt_dst_data63, sc2mac_wt_dst_data64, sc2mac_wt_dst_data65, sc2mac_wt_dst_data66, sc2mac_wt_dst_data67, sc2mac_wt_dst_data68, sc2mac_wt_dst_data69, sc2mac_wt_dst_data70, sc2mac_wt_dst_data71, sc2mac_wt_dst_data72, sc2mac_wt_dst_data73, sc2mac_wt_dst_data74, sc2mac_wt_dst_data75, sc2mac_wt_dst_data76, sc2mac_wt_dst_data77, sc2mac_wt_dst_data78, sc2mac_wt_dst_data79, sc2mac_wt_dst_data80, sc2mac_wt_dst_data81, sc2mac_wt_dst_data82, sc2mac_wt_dst_data83, sc2mac_wt_dst_data84, sc2mac_wt_dst_data85, sc2mac_wt_dst_data86, sc2mac_wt_dst_data87, sc2mac_wt_dst_data88, sc2mac_wt_dst_data89, sc2mac_wt_dst_data90, sc2mac_wt_dst_data91, sc2mac_wt_dst_data92, sc2mac_wt_dst_data93, sc2mac_wt_dst_data94, sc2mac_wt_dst_data95, sc2mac_wt_dst_data96, sc2mac_wt_dst_data97, sc2mac_wt_dst_data98, sc2mac_wt_dst_data99, sc2mac_wt_dst_data100, sc2mac_wt_dst_data101, sc2mac_wt_dst_data102, sc2mac_wt_dst_data103, sc2mac_wt_dst_data104, sc2mac_wt_dst_data105, sc2mac_wt_dst_data106, sc2mac_wt_dst_data107, sc2mac_wt_dst_data108, sc2mac_wt_dst_data109, sc2mac_wt_dst_data110, sc2mac_wt_dst_data111, sc2mac_wt_dst_data112, sc2mac_wt_dst_data113, sc2mac_wt_dst_data114, sc2mac_wt_dst_data115, sc2mac_wt_dst_data116, sc2mac_wt_dst_data117, sc2mac_wt_dst_data118, sc2mac_wt_dst_data119, sc2mac_wt_dst_data120, sc2mac_wt_dst_data121, sc2mac_wt_dst_data122, sc2mac_wt_dst_data123, sc2mac_wt_dst_data124, sc2mac_wt_dst_data125, sc2mac_wt_dst_data126, sc2mac_wt_dst_data127, sc2mac_wt_dst_sel, sc2mac_dat_dst_pvld, sc2mac_dat_dst_mask, sc2mac_dat_dst_data0, sc2mac_dat_dst_data1, sc2mac_dat_dst_data2, sc2mac_dat_dst_data3, sc2mac_dat_dst_data4, sc2mac_dat_dst_data5, sc2mac_dat_dst_data6, sc2mac_dat_dst_data7, sc2mac_dat_dst_data8, sc2mac_dat_dst_data9, sc2mac_dat_dst_data10, sc2mac_dat_dst_data11, sc2mac_dat_dst_data12, sc2mac_dat_dst_data13, sc2mac_dat_dst_data14, sc2mac_dat_dst_data15, sc2mac_dat_dst_data16, sc2mac_dat_dst_data17, sc2mac_dat_dst_data18, sc2mac_dat_dst_data19, sc2mac_dat_dst_data20, sc2mac_dat_dst_data21, sc2mac_dat_dst_data22, sc2mac_dat_dst_data23, sc2mac_dat_dst_data24, sc2mac_dat_dst_data25, sc2mac_dat_dst_data26, sc2mac_dat_dst_data27, sc2mac_dat_dst_data28, sc2mac_dat_dst_data29, sc2mac_dat_dst_data30, sc2mac_dat_dst_data31, sc2mac_dat_dst_data32, sc2mac_dat_dst_data33, sc2mac_dat_dst_data34, sc2mac_dat_dst_data35, sc2mac_dat_dst_data36, sc2mac_dat_dst_data37, sc2mac_dat_dst_data38, sc2mac_dat_dst_data39, sc2mac_dat_dst_data40, sc2mac_dat_dst_data41, sc2mac_dat_dst_data42, sc2mac_dat_dst_data43, sc2mac_dat_dst_data44, sc2mac_dat_dst_data45, sc2mac_dat_dst_data46, sc2mac_dat_dst_data47, sc2mac_dat_dst_data48, sc2mac_dat_dst_data49, sc2mac_dat_dst_data50, sc2mac_dat_dst_data51, sc2mac_dat_dst_data52, sc2mac_dat_dst_data53, sc2mac_dat_dst_data54, sc2mac_dat_dst_data55, sc2mac_dat_dst_data56, sc2mac_dat_dst_data57, sc2mac_dat_dst_data58, sc2mac_dat_dst_data59, sc2mac_dat_dst_data60, sc2mac_dat_dst_data61, sc2mac_dat_dst_data62, sc2mac_dat_dst_data63, sc2mac_dat_dst_data64, sc2mac_dat_dst_data65, sc2mac_dat_dst_data66, sc2mac_dat_dst_data67, sc2mac_dat_dst_data68, sc2mac_dat_dst_data69, sc2mac_dat_dst_data70, sc2mac_dat_dst_data71, sc2mac_dat_dst_data72, sc2mac_dat_dst_data73, sc2mac_dat_dst_data74, sc2mac_dat_dst_data75, sc2mac_dat_dst_data76, sc2mac_dat_dst_data77, sc2mac_dat_dst_data78, sc2mac_dat_dst_data79, sc2mac_dat_dst_data80, sc2mac_dat_dst_data81, sc2mac_dat_dst_data82, sc2mac_dat_dst_data83, sc2mac_dat_dst_data84, sc2mac_dat_dst_data85, sc2mac_dat_dst_data86, sc2mac_dat_dst_data87, sc2mac_dat_dst_data88, sc2mac_dat_dst_data89, sc2mac_dat_dst_data90, sc2mac_dat_dst_data91, sc2mac_dat_dst_data92, sc2mac_dat_dst_data93, sc2mac_dat_dst_data94, sc2mac_dat_dst_data95, sc2mac_dat_dst_data96, sc2mac_dat_dst_data97, sc2mac_dat_dst_data98, sc2mac_dat_dst_data99, sc2mac_dat_dst_data100, sc2mac_dat_dst_data101, sc2mac_dat_dst_data102, sc2mac_dat_dst_data103, sc2mac_dat_dst_data104, sc2mac_dat_dst_data105, sc2mac_dat_dst_data106, sc2mac_dat_dst_data107, sc2mac_dat_dst_data108, sc2mac_dat_dst_data109, sc2mac_dat_dst_data110, sc2mac_dat_dst_data111, sc2mac_dat_dst_data112, sc2mac_dat_dst_data113, sc2mac_dat_dst_data114, sc2mac_dat_dst_data115, sc2mac_dat_dst_data116, sc2mac_dat_dst_data117, sc2mac_dat_dst_data118, sc2mac_dat_dst_data119, sc2mac_dat_dst_data120, sc2mac_dat_dst_data121, sc2mac_dat_dst_data122, sc2mac_dat_dst_data123, sc2mac_dat_dst_data124, sc2mac_dat_dst_data125, sc2mac_dat_dst_data126, sc2mac_dat_dst_data127, sc2mac_dat_dst_pd);
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3390" *)
  wire [7:0] _000_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4390" *)
  wire [7:0] _001_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4400" *)
  wire [7:0] _002_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4410" *)
  wire [7:0] _003_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4420" *)
  wire [7:0] _004_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4430" *)
  wire [7:0] _005_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4440" *)
  wire [7:0] _006_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4450" *)
  wire [7:0] _007_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4460" *)
  wire [7:0] _008_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4470" *)
  wire [7:0] _009_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4480" *)
  wire [7:0] _010_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3490" *)
  wire [7:0] _011_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4490" *)
  wire [7:0] _012_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4500" *)
  wire [7:0] _013_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4510" *)
  wire [7:0] _014_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4520" *)
  wire [7:0] _015_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4530" *)
  wire [7:0] _016_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4540" *)
  wire [7:0] _017_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4550" *)
  wire [7:0] _018_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4560" *)
  wire [7:0] _019_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4570" *)
  wire [7:0] _020_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4580" *)
  wire [7:0] _021_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3500" *)
  wire [7:0] _022_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4590" *)
  wire [7:0] _023_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4600" *)
  wire [7:0] _024_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4610" *)
  wire [7:0] _025_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4620" *)
  wire [7:0] _026_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4630" *)
  wire [7:0] _027_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4640" *)
  wire [7:0] _028_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4650" *)
  wire [7:0] _029_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4660" *)
  wire [7:0] _030_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3510" *)
  wire [7:0] _031_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3520" *)
  wire [7:0] _032_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3530" *)
  wire [7:0] _033_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3540" *)
  wire [7:0] _034_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3550" *)
  wire [7:0] _035_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3560" *)
  wire [7:0] _036_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3570" *)
  wire [7:0] _037_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3580" *)
  wire [7:0] _038_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3400" *)
  wire [7:0] _039_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3590" *)
  wire [7:0] _040_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3600" *)
  wire [7:0] _041_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3610" *)
  wire [7:0] _042_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3620" *)
  wire [7:0] _043_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3630" *)
  wire [7:0] _044_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3640" *)
  wire [7:0] _045_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3650" *)
  wire [7:0] _046_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3660" *)
  wire [7:0] _047_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3670" *)
  wire [7:0] _048_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3680" *)
  wire [7:0] _049_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3410" *)
  wire [7:0] _050_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3690" *)
  wire [7:0] _051_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3700" *)
  wire [7:0] _052_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3710" *)
  wire [7:0] _053_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3720" *)
  wire [7:0] _054_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3730" *)
  wire [7:0] _055_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3740" *)
  wire [7:0] _056_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3750" *)
  wire [7:0] _057_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3760" *)
  wire [7:0] _058_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3770" *)
  wire [7:0] _059_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3780" *)
  wire [7:0] _060_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3420" *)
  wire [7:0] _061_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3790" *)
  wire [7:0] _062_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3800" *)
  wire [7:0] _063_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3810" *)
  wire [7:0] _064_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3820" *)
  wire [7:0] _065_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3830" *)
  wire [7:0] _066_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3840" *)
  wire [7:0] _067_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3850" *)
  wire [7:0] _068_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3860" *)
  wire [7:0] _069_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3870" *)
  wire [7:0] _070_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3880" *)
  wire [7:0] _071_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3430" *)
  wire [7:0] _072_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3890" *)
  wire [7:0] _073_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3900" *)
  wire [7:0] _074_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3910" *)
  wire [7:0] _075_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3920" *)
  wire [7:0] _076_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3930" *)
  wire [7:0] _077_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3940" *)
  wire [7:0] _078_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3950" *)
  wire [7:0] _079_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3960" *)
  wire [7:0] _080_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3970" *)
  wire [7:0] _081_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3980" *)
  wire [7:0] _082_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3440" *)
  wire [7:0] _083_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3990" *)
  wire [7:0] _084_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4000" *)
  wire [7:0] _085_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4010" *)
  wire [7:0] _086_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4020" *)
  wire [7:0] _087_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4030" *)
  wire [7:0] _088_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4040" *)
  wire [7:0] _089_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4050" *)
  wire [7:0] _090_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4060" *)
  wire [7:0] _091_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4070" *)
  wire [7:0] _092_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4080" *)
  wire [7:0] _093_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3450" *)
  wire [7:0] _094_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4090" *)
  wire [7:0] _095_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4100" *)
  wire [7:0] _096_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4110" *)
  wire [7:0] _097_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4120" *)
  wire [7:0] _098_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4130" *)
  wire [7:0] _099_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4140" *)
  wire [7:0] _100_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4150" *)
  wire [7:0] _101_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4160" *)
  wire [7:0] _102_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4170" *)
  wire [7:0] _103_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4180" *)
  wire [7:0] _104_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3460" *)
  wire [7:0] _105_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4190" *)
  wire [7:0] _106_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4200" *)
  wire [7:0] _107_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4210" *)
  wire [7:0] _108_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4220" *)
  wire [7:0] _109_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4230" *)
  wire [7:0] _110_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4240" *)
  wire [7:0] _111_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4250" *)
  wire [7:0] _112_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4260" *)
  wire [7:0] _113_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4270" *)
  wire [7:0] _114_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4280" *)
  wire [7:0] _115_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3470" *)
  wire [7:0] _116_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4290" *)
  wire [7:0] _117_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4300" *)
  wire [7:0] _118_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4310" *)
  wire [7:0] _119_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4320" *)
  wire [7:0] _120_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4330" *)
  wire [7:0] _121_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4340" *)
  wire [7:0] _122_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4350" *)
  wire [7:0] _123_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4360" *)
  wire [7:0] _124_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4370" *)
  wire [7:0] _125_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4380" *)
  wire [7:0] _126_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3480" *)
  wire [7:0] _127_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3329" *)
  wire [127:0] _128_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3268" *)
  wire [8:0] _129_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1981" *)
  wire [7:0] _130_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2981" *)
  wire [7:0] _131_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2991" *)
  wire [7:0] _132_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3001" *)
  wire [7:0] _133_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3011" *)
  wire [7:0] _134_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3021" *)
  wire [7:0] _135_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3031" *)
  wire [7:0] _136_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3041" *)
  wire [7:0] _137_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3051" *)
  wire [7:0] _138_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3061" *)
  wire [7:0] _139_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3071" *)
  wire [7:0] _140_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2081" *)
  wire [7:0] _141_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3081" *)
  wire [7:0] _142_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3091" *)
  wire [7:0] _143_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3101" *)
  wire [7:0] _144_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3111" *)
  wire [7:0] _145_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3121" *)
  wire [7:0] _146_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3131" *)
  wire [7:0] _147_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3141" *)
  wire [7:0] _148_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3151" *)
  wire [7:0] _149_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3161" *)
  wire [7:0] _150_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3171" *)
  wire [7:0] _151_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2091" *)
  wire [7:0] _152_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3181" *)
  wire [7:0] _153_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3191" *)
  wire [7:0] _154_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3201" *)
  wire [7:0] _155_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3211" *)
  wire [7:0] _156_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3221" *)
  wire [7:0] _157_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3231" *)
  wire [7:0] _158_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3241" *)
  wire [7:0] _159_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3251" *)
  wire [7:0] _160_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2101" *)
  wire [7:0] _161_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2111" *)
  wire [7:0] _162_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2121" *)
  wire [7:0] _163_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2131" *)
  wire [7:0] _164_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2141" *)
  wire [7:0] _165_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2151" *)
  wire [7:0] _166_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2161" *)
  wire [7:0] _167_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2171" *)
  wire [7:0] _168_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1991" *)
  wire [7:0] _169_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2181" *)
  wire [7:0] _170_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2191" *)
  wire [7:0] _171_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2201" *)
  wire [7:0] _172_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2211" *)
  wire [7:0] _173_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2221" *)
  wire [7:0] _174_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2231" *)
  wire [7:0] _175_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2241" *)
  wire [7:0] _176_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2251" *)
  wire [7:0] _177_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2261" *)
  wire [7:0] _178_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2271" *)
  wire [7:0] _179_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2001" *)
  wire [7:0] _180_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2281" *)
  wire [7:0] _181_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2291" *)
  wire [7:0] _182_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2301" *)
  wire [7:0] _183_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2311" *)
  wire [7:0] _184_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2321" *)
  wire [7:0] _185_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2331" *)
  wire [7:0] _186_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2341" *)
  wire [7:0] _187_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2351" *)
  wire [7:0] _188_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2361" *)
  wire [7:0] _189_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2371" *)
  wire [7:0] _190_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2011" *)
  wire [7:0] _191_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2381" *)
  wire [7:0] _192_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2391" *)
  wire [7:0] _193_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2401" *)
  wire [7:0] _194_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2411" *)
  wire [7:0] _195_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2421" *)
  wire [7:0] _196_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2431" *)
  wire [7:0] _197_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2441" *)
  wire [7:0] _198_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2451" *)
  wire [7:0] _199_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2461" *)
  wire [7:0] _200_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2471" *)
  wire [7:0] _201_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2021" *)
  wire [7:0] _202_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2481" *)
  wire [7:0] _203_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2491" *)
  wire [7:0] _204_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2501" *)
  wire [7:0] _205_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2511" *)
  wire [7:0] _206_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2521" *)
  wire [7:0] _207_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2531" *)
  wire [7:0] _208_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2541" *)
  wire [7:0] _209_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2551" *)
  wire [7:0] _210_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2561" *)
  wire [7:0] _211_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2571" *)
  wire [7:0] _212_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2031" *)
  wire [7:0] _213_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2581" *)
  wire [7:0] _214_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2591" *)
  wire [7:0] _215_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2601" *)
  wire [7:0] _216_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2611" *)
  wire [7:0] _217_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2621" *)
  wire [7:0] _218_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2631" *)
  wire [7:0] _219_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2641" *)
  wire [7:0] _220_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2651" *)
  wire [7:0] _221_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2661" *)
  wire [7:0] _222_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2671" *)
  wire [7:0] _223_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2041" *)
  wire [7:0] _224_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2681" *)
  wire [7:0] _225_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2691" *)
  wire [7:0] _226_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2701" *)
  wire [7:0] _227_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2711" *)
  wire [7:0] _228_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2721" *)
  wire [7:0] _229_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2731" *)
  wire [7:0] _230_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2741" *)
  wire [7:0] _231_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2751" *)
  wire [7:0] _232_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2761" *)
  wire [7:0] _233_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2771" *)
  wire [7:0] _234_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2051" *)
  wire [7:0] _235_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2781" *)
  wire [7:0] _236_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2791" *)
  wire [7:0] _237_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2801" *)
  wire [7:0] _238_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2811" *)
  wire [7:0] _239_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2821" *)
  wire [7:0] _240_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2831" *)
  wire [7:0] _241_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2841" *)
  wire [7:0] _242_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2851" *)
  wire [7:0] _243_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2861" *)
  wire [7:0] _244_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2871" *)
  wire [7:0] _245_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2061" *)
  wire [7:0] _246_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2881" *)
  wire [7:0] _247_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2891" *)
  wire [7:0] _248_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2901" *)
  wire [7:0] _249_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2911" *)
  wire [7:0] _250_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2921" *)
  wire [7:0] _251_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2931" *)
  wire [7:0] _252_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2941" *)
  wire [7:0] _253_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2951" *)
  wire [7:0] _254_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2961" *)
  wire [7:0] _255_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2971" *)
  wire [7:0] _256_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2071" *)
  wire [7:0] _257_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1920" *)
  wire [127:0] _258_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1859" *)
  wire [7:0] _259_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1863" *)
  wire _260_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3272" *)
  wire _261_;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:540" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:541" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1066" *)
  wire [7:0] sc2mac_dat_data0_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1328" *)
  reg [7:0] sc2mac_dat_data0_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1067" *)
  wire [7:0] sc2mac_dat_data100_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1329" *)
  reg [7:0] sc2mac_dat_data100_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1068" *)
  wire [7:0] sc2mac_dat_data101_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1330" *)
  reg [7:0] sc2mac_dat_data101_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1069" *)
  wire [7:0] sc2mac_dat_data102_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1331" *)
  reg [7:0] sc2mac_dat_data102_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1070" *)
  wire [7:0] sc2mac_dat_data103_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1332" *)
  reg [7:0] sc2mac_dat_data103_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1071" *)
  wire [7:0] sc2mac_dat_data104_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1333" *)
  reg [7:0] sc2mac_dat_data104_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1072" *)
  wire [7:0] sc2mac_dat_data105_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1334" *)
  reg [7:0] sc2mac_dat_data105_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1073" *)
  wire [7:0] sc2mac_dat_data106_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1335" *)
  reg [7:0] sc2mac_dat_data106_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1074" *)
  wire [7:0] sc2mac_dat_data107_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1336" *)
  reg [7:0] sc2mac_dat_data107_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1075" *)
  wire [7:0] sc2mac_dat_data108_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1337" *)
  reg [7:0] sc2mac_dat_data108_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1076" *)
  wire [7:0] sc2mac_dat_data109_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1338" *)
  reg [7:0] sc2mac_dat_data109_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1077" *)
  wire [7:0] sc2mac_dat_data10_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1339" *)
  reg [7:0] sc2mac_dat_data10_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1078" *)
  wire [7:0] sc2mac_dat_data110_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1340" *)
  reg [7:0] sc2mac_dat_data110_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1079" *)
  wire [7:0] sc2mac_dat_data111_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1341" *)
  reg [7:0] sc2mac_dat_data111_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1080" *)
  wire [7:0] sc2mac_dat_data112_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1342" *)
  reg [7:0] sc2mac_dat_data112_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1081" *)
  wire [7:0] sc2mac_dat_data113_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1343" *)
  reg [7:0] sc2mac_dat_data113_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1082" *)
  wire [7:0] sc2mac_dat_data114_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1344" *)
  reg [7:0] sc2mac_dat_data114_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1083" *)
  wire [7:0] sc2mac_dat_data115_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1345" *)
  reg [7:0] sc2mac_dat_data115_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1084" *)
  wire [7:0] sc2mac_dat_data116_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1346" *)
  reg [7:0] sc2mac_dat_data116_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1085" *)
  wire [7:0] sc2mac_dat_data117_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1347" *)
  reg [7:0] sc2mac_dat_data117_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1086" *)
  wire [7:0] sc2mac_dat_data118_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1348" *)
  reg [7:0] sc2mac_dat_data118_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1087" *)
  wire [7:0] sc2mac_dat_data119_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1349" *)
  reg [7:0] sc2mac_dat_data119_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1088" *)
  wire [7:0] sc2mac_dat_data11_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1350" *)
  reg [7:0] sc2mac_dat_data11_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1089" *)
  wire [7:0] sc2mac_dat_data120_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1351" *)
  reg [7:0] sc2mac_dat_data120_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1090" *)
  wire [7:0] sc2mac_dat_data121_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1352" *)
  reg [7:0] sc2mac_dat_data121_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1091" *)
  wire [7:0] sc2mac_dat_data122_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1353" *)
  reg [7:0] sc2mac_dat_data122_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1092" *)
  wire [7:0] sc2mac_dat_data123_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1354" *)
  reg [7:0] sc2mac_dat_data123_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1093" *)
  wire [7:0] sc2mac_dat_data124_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1355" *)
  reg [7:0] sc2mac_dat_data124_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1094" *)
  wire [7:0] sc2mac_dat_data125_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1356" *)
  reg [7:0] sc2mac_dat_data125_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1095" *)
  wire [7:0] sc2mac_dat_data126_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1357" *)
  reg [7:0] sc2mac_dat_data126_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1096" *)
  wire [7:0] sc2mac_dat_data127_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1358" *)
  reg [7:0] sc2mac_dat_data127_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1097" *)
  wire [7:0] sc2mac_dat_data12_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1359" *)
  reg [7:0] sc2mac_dat_data12_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1098" *)
  wire [7:0] sc2mac_dat_data13_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1360" *)
  reg [7:0] sc2mac_dat_data13_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1099" *)
  wire [7:0] sc2mac_dat_data14_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1361" *)
  reg [7:0] sc2mac_dat_data14_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1100" *)
  wire [7:0] sc2mac_dat_data15_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1362" *)
  reg [7:0] sc2mac_dat_data15_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1101" *)
  wire [7:0] sc2mac_dat_data16_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1363" *)
  reg [7:0] sc2mac_dat_data16_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1102" *)
  wire [7:0] sc2mac_dat_data17_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1364" *)
  reg [7:0] sc2mac_dat_data17_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1103" *)
  wire [7:0] sc2mac_dat_data18_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1365" *)
  reg [7:0] sc2mac_dat_data18_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1104" *)
  wire [7:0] sc2mac_dat_data19_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1366" *)
  reg [7:0] sc2mac_dat_data19_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1105" *)
  wire [7:0] sc2mac_dat_data1_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1367" *)
  reg [7:0] sc2mac_dat_data1_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1106" *)
  wire [7:0] sc2mac_dat_data20_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1368" *)
  reg [7:0] sc2mac_dat_data20_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1107" *)
  wire [7:0] sc2mac_dat_data21_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1369" *)
  reg [7:0] sc2mac_dat_data21_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1108" *)
  wire [7:0] sc2mac_dat_data22_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1370" *)
  reg [7:0] sc2mac_dat_data22_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1109" *)
  wire [7:0] sc2mac_dat_data23_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1371" *)
  reg [7:0] sc2mac_dat_data23_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1110" *)
  wire [7:0] sc2mac_dat_data24_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1372" *)
  reg [7:0] sc2mac_dat_data24_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1111" *)
  wire [7:0] sc2mac_dat_data25_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1373" *)
  reg [7:0] sc2mac_dat_data25_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1112" *)
  wire [7:0] sc2mac_dat_data26_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1374" *)
  reg [7:0] sc2mac_dat_data26_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1113" *)
  wire [7:0] sc2mac_dat_data27_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1375" *)
  reg [7:0] sc2mac_dat_data27_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1114" *)
  wire [7:0] sc2mac_dat_data28_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1376" *)
  reg [7:0] sc2mac_dat_data28_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1115" *)
  wire [7:0] sc2mac_dat_data29_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1377" *)
  reg [7:0] sc2mac_dat_data29_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1116" *)
  wire [7:0] sc2mac_dat_data2_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1378" *)
  reg [7:0] sc2mac_dat_data2_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1117" *)
  wire [7:0] sc2mac_dat_data30_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1379" *)
  reg [7:0] sc2mac_dat_data30_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1118" *)
  wire [7:0] sc2mac_dat_data31_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1380" *)
  reg [7:0] sc2mac_dat_data31_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1119" *)
  wire [7:0] sc2mac_dat_data32_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1381" *)
  reg [7:0] sc2mac_dat_data32_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1120" *)
  wire [7:0] sc2mac_dat_data33_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1382" *)
  reg [7:0] sc2mac_dat_data33_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1121" *)
  wire [7:0] sc2mac_dat_data34_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1383" *)
  reg [7:0] sc2mac_dat_data34_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1122" *)
  wire [7:0] sc2mac_dat_data35_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1384" *)
  reg [7:0] sc2mac_dat_data35_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1123" *)
  wire [7:0] sc2mac_dat_data36_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1385" *)
  reg [7:0] sc2mac_dat_data36_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1124" *)
  wire [7:0] sc2mac_dat_data37_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1386" *)
  reg [7:0] sc2mac_dat_data37_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1125" *)
  wire [7:0] sc2mac_dat_data38_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1387" *)
  reg [7:0] sc2mac_dat_data38_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1126" *)
  wire [7:0] sc2mac_dat_data39_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1388" *)
  reg [7:0] sc2mac_dat_data39_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1127" *)
  wire [7:0] sc2mac_dat_data3_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1389" *)
  reg [7:0] sc2mac_dat_data3_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1128" *)
  wire [7:0] sc2mac_dat_data40_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1390" *)
  reg [7:0] sc2mac_dat_data40_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1129" *)
  wire [7:0] sc2mac_dat_data41_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1391" *)
  reg [7:0] sc2mac_dat_data41_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1130" *)
  wire [7:0] sc2mac_dat_data42_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1392" *)
  reg [7:0] sc2mac_dat_data42_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1131" *)
  wire [7:0] sc2mac_dat_data43_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1393" *)
  reg [7:0] sc2mac_dat_data43_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1132" *)
  wire [7:0] sc2mac_dat_data44_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1394" *)
  reg [7:0] sc2mac_dat_data44_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1133" *)
  wire [7:0] sc2mac_dat_data45_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1395" *)
  reg [7:0] sc2mac_dat_data45_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1134" *)
  wire [7:0] sc2mac_dat_data46_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1396" *)
  reg [7:0] sc2mac_dat_data46_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1135" *)
  wire [7:0] sc2mac_dat_data47_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1397" *)
  reg [7:0] sc2mac_dat_data47_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1136" *)
  wire [7:0] sc2mac_dat_data48_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1398" *)
  reg [7:0] sc2mac_dat_data48_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1137" *)
  wire [7:0] sc2mac_dat_data49_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1399" *)
  reg [7:0] sc2mac_dat_data49_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1138" *)
  wire [7:0] sc2mac_dat_data4_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1400" *)
  reg [7:0] sc2mac_dat_data4_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1139" *)
  wire [7:0] sc2mac_dat_data50_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1401" *)
  reg [7:0] sc2mac_dat_data50_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1140" *)
  wire [7:0] sc2mac_dat_data51_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1402" *)
  reg [7:0] sc2mac_dat_data51_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1141" *)
  wire [7:0] sc2mac_dat_data52_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1403" *)
  reg [7:0] sc2mac_dat_data52_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1142" *)
  wire [7:0] sc2mac_dat_data53_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1404" *)
  reg [7:0] sc2mac_dat_data53_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1143" *)
  wire [7:0] sc2mac_dat_data54_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1405" *)
  reg [7:0] sc2mac_dat_data54_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1144" *)
  wire [7:0] sc2mac_dat_data55_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1406" *)
  reg [7:0] sc2mac_dat_data55_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1145" *)
  wire [7:0] sc2mac_dat_data56_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1407" *)
  reg [7:0] sc2mac_dat_data56_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1146" *)
  wire [7:0] sc2mac_dat_data57_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1408" *)
  reg [7:0] sc2mac_dat_data57_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1147" *)
  wire [7:0] sc2mac_dat_data58_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1409" *)
  reg [7:0] sc2mac_dat_data58_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1148" *)
  wire [7:0] sc2mac_dat_data59_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1410" *)
  reg [7:0] sc2mac_dat_data59_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1149" *)
  wire [7:0] sc2mac_dat_data5_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1411" *)
  reg [7:0] sc2mac_dat_data5_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1150" *)
  wire [7:0] sc2mac_dat_data60_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1412" *)
  reg [7:0] sc2mac_dat_data60_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1151" *)
  wire [7:0] sc2mac_dat_data61_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1413" *)
  reg [7:0] sc2mac_dat_data61_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1152" *)
  wire [7:0] sc2mac_dat_data62_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1414" *)
  reg [7:0] sc2mac_dat_data62_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1153" *)
  wire [7:0] sc2mac_dat_data63_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1415" *)
  reg [7:0] sc2mac_dat_data63_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1154" *)
  wire [7:0] sc2mac_dat_data64_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1416" *)
  reg [7:0] sc2mac_dat_data64_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1155" *)
  wire [7:0] sc2mac_dat_data65_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1417" *)
  reg [7:0] sc2mac_dat_data65_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1156" *)
  wire [7:0] sc2mac_dat_data66_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1418" *)
  reg [7:0] sc2mac_dat_data66_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1157" *)
  wire [7:0] sc2mac_dat_data67_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1419" *)
  reg [7:0] sc2mac_dat_data67_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1158" *)
  wire [7:0] sc2mac_dat_data68_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1420" *)
  reg [7:0] sc2mac_dat_data68_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1159" *)
  wire [7:0] sc2mac_dat_data69_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1421" *)
  reg [7:0] sc2mac_dat_data69_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1160" *)
  wire [7:0] sc2mac_dat_data6_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1422" *)
  reg [7:0] sc2mac_dat_data6_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1161" *)
  wire [7:0] sc2mac_dat_data70_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1423" *)
  reg [7:0] sc2mac_dat_data70_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1162" *)
  wire [7:0] sc2mac_dat_data71_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1424" *)
  reg [7:0] sc2mac_dat_data71_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1163" *)
  wire [7:0] sc2mac_dat_data72_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1425" *)
  reg [7:0] sc2mac_dat_data72_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1164" *)
  wire [7:0] sc2mac_dat_data73_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1426" *)
  reg [7:0] sc2mac_dat_data73_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1165" *)
  wire [7:0] sc2mac_dat_data74_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1427" *)
  reg [7:0] sc2mac_dat_data74_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1166" *)
  wire [7:0] sc2mac_dat_data75_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1428" *)
  reg [7:0] sc2mac_dat_data75_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1167" *)
  wire [7:0] sc2mac_dat_data76_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1429" *)
  reg [7:0] sc2mac_dat_data76_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1168" *)
  wire [7:0] sc2mac_dat_data77_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1430" *)
  reg [7:0] sc2mac_dat_data77_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1169" *)
  wire [7:0] sc2mac_dat_data78_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1431" *)
  reg [7:0] sc2mac_dat_data78_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1170" *)
  wire [7:0] sc2mac_dat_data79_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1432" *)
  reg [7:0] sc2mac_dat_data79_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1171" *)
  wire [7:0] sc2mac_dat_data7_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1433" *)
  reg [7:0] sc2mac_dat_data7_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1172" *)
  wire [7:0] sc2mac_dat_data80_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1434" *)
  reg [7:0] sc2mac_dat_data80_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1173" *)
  wire [7:0] sc2mac_dat_data81_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1435" *)
  reg [7:0] sc2mac_dat_data81_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1174" *)
  wire [7:0] sc2mac_dat_data82_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1436" *)
  reg [7:0] sc2mac_dat_data82_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1175" *)
  wire [7:0] sc2mac_dat_data83_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1437" *)
  reg [7:0] sc2mac_dat_data83_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1176" *)
  wire [7:0] sc2mac_dat_data84_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1438" *)
  reg [7:0] sc2mac_dat_data84_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1177" *)
  wire [7:0] sc2mac_dat_data85_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1439" *)
  reg [7:0] sc2mac_dat_data85_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1178" *)
  wire [7:0] sc2mac_dat_data86_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1440" *)
  reg [7:0] sc2mac_dat_data86_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1179" *)
  wire [7:0] sc2mac_dat_data87_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1441" *)
  reg [7:0] sc2mac_dat_data87_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1180" *)
  wire [7:0] sc2mac_dat_data88_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1442" *)
  reg [7:0] sc2mac_dat_data88_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1181" *)
  wire [7:0] sc2mac_dat_data89_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1443" *)
  reg [7:0] sc2mac_dat_data89_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1182" *)
  wire [7:0] sc2mac_dat_data8_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1444" *)
  reg [7:0] sc2mac_dat_data8_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1183" *)
  wire [7:0] sc2mac_dat_data90_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1445" *)
  reg [7:0] sc2mac_dat_data90_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1184" *)
  wire [7:0] sc2mac_dat_data91_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1446" *)
  reg [7:0] sc2mac_dat_data91_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1185" *)
  wire [7:0] sc2mac_dat_data92_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1447" *)
  reg [7:0] sc2mac_dat_data92_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1186" *)
  wire [7:0] sc2mac_dat_data93_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1448" *)
  reg [7:0] sc2mac_dat_data93_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1187" *)
  wire [7:0] sc2mac_dat_data94_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1449" *)
  reg [7:0] sc2mac_dat_data94_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1188" *)
  wire [7:0] sc2mac_dat_data95_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1450" *)
  reg [7:0] sc2mac_dat_data95_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1189" *)
  wire [7:0] sc2mac_dat_data96_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1451" *)
  reg [7:0] sc2mac_dat_data96_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1190" *)
  wire [7:0] sc2mac_dat_data97_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1452" *)
  reg [7:0] sc2mac_dat_data97_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1191" *)
  wire [7:0] sc2mac_dat_data98_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1453" *)
  reg [7:0] sc2mac_dat_data98_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1192" *)
  wire [7:0] sc2mac_dat_data99_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1454" *)
  reg [7:0] sc2mac_dat_data99_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1193" *)
  wire [7:0] sc2mac_dat_data9_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1455" *)
  reg [7:0] sc2mac_dat_data9_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:937" *)
  output [7:0] sc2mac_dat_dst_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:938" *)
  output [7:0] sc2mac_dat_dst_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:947" *)
  output [7:0] sc2mac_dat_dst_data10;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1037" *)
  output [7:0] sc2mac_dat_dst_data100;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1038" *)
  output [7:0] sc2mac_dat_dst_data101;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1039" *)
  output [7:0] sc2mac_dat_dst_data102;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1040" *)
  output [7:0] sc2mac_dat_dst_data103;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1041" *)
  output [7:0] sc2mac_dat_dst_data104;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1042" *)
  output [7:0] sc2mac_dat_dst_data105;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1043" *)
  output [7:0] sc2mac_dat_dst_data106;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1044" *)
  output [7:0] sc2mac_dat_dst_data107;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1045" *)
  output [7:0] sc2mac_dat_dst_data108;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1046" *)
  output [7:0] sc2mac_dat_dst_data109;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:948" *)
  output [7:0] sc2mac_dat_dst_data11;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1047" *)
  output [7:0] sc2mac_dat_dst_data110;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1048" *)
  output [7:0] sc2mac_dat_dst_data111;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1049" *)
  output [7:0] sc2mac_dat_dst_data112;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1050" *)
  output [7:0] sc2mac_dat_dst_data113;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1051" *)
  output [7:0] sc2mac_dat_dst_data114;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1052" *)
  output [7:0] sc2mac_dat_dst_data115;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1053" *)
  output [7:0] sc2mac_dat_dst_data116;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1054" *)
  output [7:0] sc2mac_dat_dst_data117;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1055" *)
  output [7:0] sc2mac_dat_dst_data118;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1056" *)
  output [7:0] sc2mac_dat_dst_data119;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:949" *)
  output [7:0] sc2mac_dat_dst_data12;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1057" *)
  output [7:0] sc2mac_dat_dst_data120;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1058" *)
  output [7:0] sc2mac_dat_dst_data121;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1059" *)
  output [7:0] sc2mac_dat_dst_data122;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1060" *)
  output [7:0] sc2mac_dat_dst_data123;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1061" *)
  output [7:0] sc2mac_dat_dst_data124;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1062" *)
  output [7:0] sc2mac_dat_dst_data125;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1063" *)
  output [7:0] sc2mac_dat_dst_data126;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1064" *)
  output [7:0] sc2mac_dat_dst_data127;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:950" *)
  output [7:0] sc2mac_dat_dst_data13;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:951" *)
  output [7:0] sc2mac_dat_dst_data14;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:952" *)
  output [7:0] sc2mac_dat_dst_data15;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:953" *)
  output [7:0] sc2mac_dat_dst_data16;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:954" *)
  output [7:0] sc2mac_dat_dst_data17;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:955" *)
  output [7:0] sc2mac_dat_dst_data18;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:956" *)
  output [7:0] sc2mac_dat_dst_data19;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:939" *)
  output [7:0] sc2mac_dat_dst_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:957" *)
  output [7:0] sc2mac_dat_dst_data20;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:958" *)
  output [7:0] sc2mac_dat_dst_data21;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:959" *)
  output [7:0] sc2mac_dat_dst_data22;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:960" *)
  output [7:0] sc2mac_dat_dst_data23;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:961" *)
  output [7:0] sc2mac_dat_dst_data24;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:962" *)
  output [7:0] sc2mac_dat_dst_data25;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:963" *)
  output [7:0] sc2mac_dat_dst_data26;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:964" *)
  output [7:0] sc2mac_dat_dst_data27;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:965" *)
  output [7:0] sc2mac_dat_dst_data28;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:966" *)
  output [7:0] sc2mac_dat_dst_data29;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:940" *)
  output [7:0] sc2mac_dat_dst_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:967" *)
  output [7:0] sc2mac_dat_dst_data30;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:968" *)
  output [7:0] sc2mac_dat_dst_data31;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:969" *)
  output [7:0] sc2mac_dat_dst_data32;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:970" *)
  output [7:0] sc2mac_dat_dst_data33;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:971" *)
  output [7:0] sc2mac_dat_dst_data34;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:972" *)
  output [7:0] sc2mac_dat_dst_data35;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:973" *)
  output [7:0] sc2mac_dat_dst_data36;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:974" *)
  output [7:0] sc2mac_dat_dst_data37;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:975" *)
  output [7:0] sc2mac_dat_dst_data38;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:976" *)
  output [7:0] sc2mac_dat_dst_data39;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:941" *)
  output [7:0] sc2mac_dat_dst_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:977" *)
  output [7:0] sc2mac_dat_dst_data40;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:978" *)
  output [7:0] sc2mac_dat_dst_data41;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:979" *)
  output [7:0] sc2mac_dat_dst_data42;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:980" *)
  output [7:0] sc2mac_dat_dst_data43;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:981" *)
  output [7:0] sc2mac_dat_dst_data44;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:982" *)
  output [7:0] sc2mac_dat_dst_data45;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:983" *)
  output [7:0] sc2mac_dat_dst_data46;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:984" *)
  output [7:0] sc2mac_dat_dst_data47;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:985" *)
  output [7:0] sc2mac_dat_dst_data48;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:986" *)
  output [7:0] sc2mac_dat_dst_data49;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:942" *)
  output [7:0] sc2mac_dat_dst_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:987" *)
  output [7:0] sc2mac_dat_dst_data50;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:988" *)
  output [7:0] sc2mac_dat_dst_data51;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:989" *)
  output [7:0] sc2mac_dat_dst_data52;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:990" *)
  output [7:0] sc2mac_dat_dst_data53;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:991" *)
  output [7:0] sc2mac_dat_dst_data54;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:992" *)
  output [7:0] sc2mac_dat_dst_data55;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:993" *)
  output [7:0] sc2mac_dat_dst_data56;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:994" *)
  output [7:0] sc2mac_dat_dst_data57;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:995" *)
  output [7:0] sc2mac_dat_dst_data58;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:996" *)
  output [7:0] sc2mac_dat_dst_data59;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:943" *)
  output [7:0] sc2mac_dat_dst_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:997" *)
  output [7:0] sc2mac_dat_dst_data60;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:998" *)
  output [7:0] sc2mac_dat_dst_data61;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:999" *)
  output [7:0] sc2mac_dat_dst_data62;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1000" *)
  output [7:0] sc2mac_dat_dst_data63;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1001" *)
  output [7:0] sc2mac_dat_dst_data64;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1002" *)
  output [7:0] sc2mac_dat_dst_data65;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1003" *)
  output [7:0] sc2mac_dat_dst_data66;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1004" *)
  output [7:0] sc2mac_dat_dst_data67;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1005" *)
  output [7:0] sc2mac_dat_dst_data68;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1006" *)
  output [7:0] sc2mac_dat_dst_data69;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:944" *)
  output [7:0] sc2mac_dat_dst_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1007" *)
  output [7:0] sc2mac_dat_dst_data70;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1008" *)
  output [7:0] sc2mac_dat_dst_data71;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1009" *)
  output [7:0] sc2mac_dat_dst_data72;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1010" *)
  output [7:0] sc2mac_dat_dst_data73;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1011" *)
  output [7:0] sc2mac_dat_dst_data74;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1012" *)
  output [7:0] sc2mac_dat_dst_data75;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1013" *)
  output [7:0] sc2mac_dat_dst_data76;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1014" *)
  output [7:0] sc2mac_dat_dst_data77;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1015" *)
  output [7:0] sc2mac_dat_dst_data78;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1016" *)
  output [7:0] sc2mac_dat_dst_data79;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:945" *)
  output [7:0] sc2mac_dat_dst_data8;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1017" *)
  output [7:0] sc2mac_dat_dst_data80;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1018" *)
  output [7:0] sc2mac_dat_dst_data81;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1019" *)
  output [7:0] sc2mac_dat_dst_data82;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1020" *)
  output [7:0] sc2mac_dat_dst_data83;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1021" *)
  output [7:0] sc2mac_dat_dst_data84;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1022" *)
  output [7:0] sc2mac_dat_dst_data85;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1023" *)
  output [7:0] sc2mac_dat_dst_data86;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1024" *)
  output [7:0] sc2mac_dat_dst_data87;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1025" *)
  output [7:0] sc2mac_dat_dst_data88;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1026" *)
  output [7:0] sc2mac_dat_dst_data89;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:946" *)
  output [7:0] sc2mac_dat_dst_data9;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1027" *)
  output [7:0] sc2mac_dat_dst_data90;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1028" *)
  output [7:0] sc2mac_dat_dst_data91;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1029" *)
  output [7:0] sc2mac_dat_dst_data92;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1030" *)
  output [7:0] sc2mac_dat_dst_data93;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1031" *)
  output [7:0] sc2mac_dat_dst_data94;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1032" *)
  output [7:0] sc2mac_dat_dst_data95;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1033" *)
  output [7:0] sc2mac_dat_dst_data96;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1034" *)
  output [7:0] sc2mac_dat_dst_data97;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1035" *)
  output [7:0] sc2mac_dat_dst_data98;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1036" *)
  output [7:0] sc2mac_dat_dst_data99;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:936" *)
  output [127:0] sc2mac_dat_dst_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1065" *)
  output [8:0] sc2mac_dat_dst_pd;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:935" *)
  output sc2mac_dat_dst_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1194" *)
  wire [127:0] sc2mac_dat_mask_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1456" *)
  reg [127:0] sc2mac_dat_mask_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1195" *)
  wire [8:0] sc2mac_dat_pd_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1457" *)
  reg [8:0] sc2mac_dat_pd_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1196" *)
  wire sc2mac_dat_pvld_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1458" *)
  reg sc2mac_dat_pvld_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:675" *)
  input [7:0] sc2mac_dat_src_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:676" *)
  input [7:0] sc2mac_dat_src_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:685" *)
  input [7:0] sc2mac_dat_src_data10;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:775" *)
  input [7:0] sc2mac_dat_src_data100;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:776" *)
  input [7:0] sc2mac_dat_src_data101;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:777" *)
  input [7:0] sc2mac_dat_src_data102;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:778" *)
  input [7:0] sc2mac_dat_src_data103;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:779" *)
  input [7:0] sc2mac_dat_src_data104;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:780" *)
  input [7:0] sc2mac_dat_src_data105;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:781" *)
  input [7:0] sc2mac_dat_src_data106;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:782" *)
  input [7:0] sc2mac_dat_src_data107;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:783" *)
  input [7:0] sc2mac_dat_src_data108;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:784" *)
  input [7:0] sc2mac_dat_src_data109;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:686" *)
  input [7:0] sc2mac_dat_src_data11;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:785" *)
  input [7:0] sc2mac_dat_src_data110;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:786" *)
  input [7:0] sc2mac_dat_src_data111;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:787" *)
  input [7:0] sc2mac_dat_src_data112;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:788" *)
  input [7:0] sc2mac_dat_src_data113;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:789" *)
  input [7:0] sc2mac_dat_src_data114;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:790" *)
  input [7:0] sc2mac_dat_src_data115;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:791" *)
  input [7:0] sc2mac_dat_src_data116;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:792" *)
  input [7:0] sc2mac_dat_src_data117;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:793" *)
  input [7:0] sc2mac_dat_src_data118;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:794" *)
  input [7:0] sc2mac_dat_src_data119;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:687" *)
  input [7:0] sc2mac_dat_src_data12;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:795" *)
  input [7:0] sc2mac_dat_src_data120;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:796" *)
  input [7:0] sc2mac_dat_src_data121;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:797" *)
  input [7:0] sc2mac_dat_src_data122;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:798" *)
  input [7:0] sc2mac_dat_src_data123;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:799" *)
  input [7:0] sc2mac_dat_src_data124;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:800" *)
  input [7:0] sc2mac_dat_src_data125;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:801" *)
  input [7:0] sc2mac_dat_src_data126;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:802" *)
  input [7:0] sc2mac_dat_src_data127;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:688" *)
  input [7:0] sc2mac_dat_src_data13;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:689" *)
  input [7:0] sc2mac_dat_src_data14;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:690" *)
  input [7:0] sc2mac_dat_src_data15;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:691" *)
  input [7:0] sc2mac_dat_src_data16;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:692" *)
  input [7:0] sc2mac_dat_src_data17;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:693" *)
  input [7:0] sc2mac_dat_src_data18;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:694" *)
  input [7:0] sc2mac_dat_src_data19;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:677" *)
  input [7:0] sc2mac_dat_src_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:695" *)
  input [7:0] sc2mac_dat_src_data20;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:696" *)
  input [7:0] sc2mac_dat_src_data21;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:697" *)
  input [7:0] sc2mac_dat_src_data22;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:698" *)
  input [7:0] sc2mac_dat_src_data23;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:699" *)
  input [7:0] sc2mac_dat_src_data24;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:700" *)
  input [7:0] sc2mac_dat_src_data25;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:701" *)
  input [7:0] sc2mac_dat_src_data26;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:702" *)
  input [7:0] sc2mac_dat_src_data27;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:703" *)
  input [7:0] sc2mac_dat_src_data28;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:704" *)
  input [7:0] sc2mac_dat_src_data29;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:678" *)
  input [7:0] sc2mac_dat_src_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:705" *)
  input [7:0] sc2mac_dat_src_data30;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:706" *)
  input [7:0] sc2mac_dat_src_data31;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:707" *)
  input [7:0] sc2mac_dat_src_data32;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:708" *)
  input [7:0] sc2mac_dat_src_data33;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:709" *)
  input [7:0] sc2mac_dat_src_data34;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:710" *)
  input [7:0] sc2mac_dat_src_data35;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:711" *)
  input [7:0] sc2mac_dat_src_data36;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:712" *)
  input [7:0] sc2mac_dat_src_data37;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:713" *)
  input [7:0] sc2mac_dat_src_data38;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:714" *)
  input [7:0] sc2mac_dat_src_data39;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:679" *)
  input [7:0] sc2mac_dat_src_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:715" *)
  input [7:0] sc2mac_dat_src_data40;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:716" *)
  input [7:0] sc2mac_dat_src_data41;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:717" *)
  input [7:0] sc2mac_dat_src_data42;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:718" *)
  input [7:0] sc2mac_dat_src_data43;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:719" *)
  input [7:0] sc2mac_dat_src_data44;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:720" *)
  input [7:0] sc2mac_dat_src_data45;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:721" *)
  input [7:0] sc2mac_dat_src_data46;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:722" *)
  input [7:0] sc2mac_dat_src_data47;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:723" *)
  input [7:0] sc2mac_dat_src_data48;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:724" *)
  input [7:0] sc2mac_dat_src_data49;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:680" *)
  input [7:0] sc2mac_dat_src_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:725" *)
  input [7:0] sc2mac_dat_src_data50;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:726" *)
  input [7:0] sc2mac_dat_src_data51;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:727" *)
  input [7:0] sc2mac_dat_src_data52;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:728" *)
  input [7:0] sc2mac_dat_src_data53;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:729" *)
  input [7:0] sc2mac_dat_src_data54;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:730" *)
  input [7:0] sc2mac_dat_src_data55;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:731" *)
  input [7:0] sc2mac_dat_src_data56;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:732" *)
  input [7:0] sc2mac_dat_src_data57;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:733" *)
  input [7:0] sc2mac_dat_src_data58;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:734" *)
  input [7:0] sc2mac_dat_src_data59;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:681" *)
  input [7:0] sc2mac_dat_src_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:735" *)
  input [7:0] sc2mac_dat_src_data60;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:736" *)
  input [7:0] sc2mac_dat_src_data61;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:737" *)
  input [7:0] sc2mac_dat_src_data62;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:738" *)
  input [7:0] sc2mac_dat_src_data63;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:739" *)
  input [7:0] sc2mac_dat_src_data64;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:740" *)
  input [7:0] sc2mac_dat_src_data65;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:741" *)
  input [7:0] sc2mac_dat_src_data66;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:742" *)
  input [7:0] sc2mac_dat_src_data67;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:743" *)
  input [7:0] sc2mac_dat_src_data68;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:744" *)
  input [7:0] sc2mac_dat_src_data69;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:682" *)
  input [7:0] sc2mac_dat_src_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:745" *)
  input [7:0] sc2mac_dat_src_data70;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:746" *)
  input [7:0] sc2mac_dat_src_data71;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:747" *)
  input [7:0] sc2mac_dat_src_data72;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:748" *)
  input [7:0] sc2mac_dat_src_data73;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:749" *)
  input [7:0] sc2mac_dat_src_data74;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:750" *)
  input [7:0] sc2mac_dat_src_data75;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:751" *)
  input [7:0] sc2mac_dat_src_data76;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:752" *)
  input [7:0] sc2mac_dat_src_data77;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:753" *)
  input [7:0] sc2mac_dat_src_data78;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:754" *)
  input [7:0] sc2mac_dat_src_data79;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:683" *)
  input [7:0] sc2mac_dat_src_data8;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:755" *)
  input [7:0] sc2mac_dat_src_data80;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:756" *)
  input [7:0] sc2mac_dat_src_data81;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:757" *)
  input [7:0] sc2mac_dat_src_data82;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:758" *)
  input [7:0] sc2mac_dat_src_data83;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:759" *)
  input [7:0] sc2mac_dat_src_data84;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:760" *)
  input [7:0] sc2mac_dat_src_data85;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:761" *)
  input [7:0] sc2mac_dat_src_data86;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:762" *)
  input [7:0] sc2mac_dat_src_data87;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:763" *)
  input [7:0] sc2mac_dat_src_data88;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:764" *)
  input [7:0] sc2mac_dat_src_data89;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:684" *)
  input [7:0] sc2mac_dat_src_data9;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:765" *)
  input [7:0] sc2mac_dat_src_data90;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:766" *)
  input [7:0] sc2mac_dat_src_data91;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:767" *)
  input [7:0] sc2mac_dat_src_data92;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:768" *)
  input [7:0] sc2mac_dat_src_data93;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:769" *)
  input [7:0] sc2mac_dat_src_data94;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:770" *)
  input [7:0] sc2mac_dat_src_data95;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:771" *)
  input [7:0] sc2mac_dat_src_data96;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:772" *)
  input [7:0] sc2mac_dat_src_data97;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:773" *)
  input [7:0] sc2mac_dat_src_data98;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:774" *)
  input [7:0] sc2mac_dat_src_data99;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:674" *)
  input [127:0] sc2mac_dat_src_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:803" *)
  input [8:0] sc2mac_dat_src_pd;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:673" *)
  input sc2mac_dat_src_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1197" *)
  wire [7:0] sc2mac_wt_data0_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1459" *)
  reg [7:0] sc2mac_wt_data0_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1198" *)
  wire [7:0] sc2mac_wt_data100_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1460" *)
  reg [7:0] sc2mac_wt_data100_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1199" *)
  wire [7:0] sc2mac_wt_data101_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1461" *)
  reg [7:0] sc2mac_wt_data101_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1200" *)
  wire [7:0] sc2mac_wt_data102_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1462" *)
  reg [7:0] sc2mac_wt_data102_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1201" *)
  wire [7:0] sc2mac_wt_data103_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1463" *)
  reg [7:0] sc2mac_wt_data103_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1202" *)
  wire [7:0] sc2mac_wt_data104_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1464" *)
  reg [7:0] sc2mac_wt_data104_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1203" *)
  wire [7:0] sc2mac_wt_data105_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1465" *)
  reg [7:0] sc2mac_wt_data105_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1204" *)
  wire [7:0] sc2mac_wt_data106_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1466" *)
  reg [7:0] sc2mac_wt_data106_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1205" *)
  wire [7:0] sc2mac_wt_data107_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1467" *)
  reg [7:0] sc2mac_wt_data107_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1206" *)
  wire [7:0] sc2mac_wt_data108_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1468" *)
  reg [7:0] sc2mac_wt_data108_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1207" *)
  wire [7:0] sc2mac_wt_data109_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1469" *)
  reg [7:0] sc2mac_wt_data109_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1208" *)
  wire [7:0] sc2mac_wt_data10_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1470" *)
  reg [7:0] sc2mac_wt_data10_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1209" *)
  wire [7:0] sc2mac_wt_data110_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1471" *)
  reg [7:0] sc2mac_wt_data110_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1210" *)
  wire [7:0] sc2mac_wt_data111_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1472" *)
  reg [7:0] sc2mac_wt_data111_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1211" *)
  wire [7:0] sc2mac_wt_data112_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1473" *)
  reg [7:0] sc2mac_wt_data112_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1212" *)
  wire [7:0] sc2mac_wt_data113_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1474" *)
  reg [7:0] sc2mac_wt_data113_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1213" *)
  wire [7:0] sc2mac_wt_data114_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1475" *)
  reg [7:0] sc2mac_wt_data114_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1214" *)
  wire [7:0] sc2mac_wt_data115_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1476" *)
  reg [7:0] sc2mac_wt_data115_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1215" *)
  wire [7:0] sc2mac_wt_data116_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1477" *)
  reg [7:0] sc2mac_wt_data116_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1216" *)
  wire [7:0] sc2mac_wt_data117_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1478" *)
  reg [7:0] sc2mac_wt_data117_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1217" *)
  wire [7:0] sc2mac_wt_data118_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1479" *)
  reg [7:0] sc2mac_wt_data118_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1218" *)
  wire [7:0] sc2mac_wt_data119_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1480" *)
  reg [7:0] sc2mac_wt_data119_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1219" *)
  wire [7:0] sc2mac_wt_data11_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1481" *)
  reg [7:0] sc2mac_wt_data11_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1220" *)
  wire [7:0] sc2mac_wt_data120_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1482" *)
  reg [7:0] sc2mac_wt_data120_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1221" *)
  wire [7:0] sc2mac_wt_data121_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1483" *)
  reg [7:0] sc2mac_wt_data121_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1222" *)
  wire [7:0] sc2mac_wt_data122_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1484" *)
  reg [7:0] sc2mac_wt_data122_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1223" *)
  wire [7:0] sc2mac_wt_data123_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1485" *)
  reg [7:0] sc2mac_wt_data123_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1224" *)
  wire [7:0] sc2mac_wt_data124_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1486" *)
  reg [7:0] sc2mac_wt_data124_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1225" *)
  wire [7:0] sc2mac_wt_data125_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1487" *)
  reg [7:0] sc2mac_wt_data125_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1226" *)
  wire [7:0] sc2mac_wt_data126_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1488" *)
  reg [7:0] sc2mac_wt_data126_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1227" *)
  wire [7:0] sc2mac_wt_data127_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1489" *)
  reg [7:0] sc2mac_wt_data127_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1228" *)
  wire [7:0] sc2mac_wt_data12_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1490" *)
  reg [7:0] sc2mac_wt_data12_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1229" *)
  wire [7:0] sc2mac_wt_data13_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1491" *)
  reg [7:0] sc2mac_wt_data13_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1230" *)
  wire [7:0] sc2mac_wt_data14_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1492" *)
  reg [7:0] sc2mac_wt_data14_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1231" *)
  wire [7:0] sc2mac_wt_data15_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1493" *)
  reg [7:0] sc2mac_wt_data15_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1232" *)
  wire [7:0] sc2mac_wt_data16_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1494" *)
  reg [7:0] sc2mac_wt_data16_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1233" *)
  wire [7:0] sc2mac_wt_data17_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1495" *)
  reg [7:0] sc2mac_wt_data17_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1234" *)
  wire [7:0] sc2mac_wt_data18_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1496" *)
  reg [7:0] sc2mac_wt_data18_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1235" *)
  wire [7:0] sc2mac_wt_data19_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1497" *)
  reg [7:0] sc2mac_wt_data19_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1236" *)
  wire [7:0] sc2mac_wt_data1_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1498" *)
  reg [7:0] sc2mac_wt_data1_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1237" *)
  wire [7:0] sc2mac_wt_data20_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1499" *)
  reg [7:0] sc2mac_wt_data20_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1238" *)
  wire [7:0] sc2mac_wt_data21_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1500" *)
  reg [7:0] sc2mac_wt_data21_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1239" *)
  wire [7:0] sc2mac_wt_data22_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1501" *)
  reg [7:0] sc2mac_wt_data22_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1240" *)
  wire [7:0] sc2mac_wt_data23_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1502" *)
  reg [7:0] sc2mac_wt_data23_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1241" *)
  wire [7:0] sc2mac_wt_data24_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1503" *)
  reg [7:0] sc2mac_wt_data24_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1242" *)
  wire [7:0] sc2mac_wt_data25_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1504" *)
  reg [7:0] sc2mac_wt_data25_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1243" *)
  wire [7:0] sc2mac_wt_data26_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1505" *)
  reg [7:0] sc2mac_wt_data26_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1244" *)
  wire [7:0] sc2mac_wt_data27_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1506" *)
  reg [7:0] sc2mac_wt_data27_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1245" *)
  wire [7:0] sc2mac_wt_data28_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1507" *)
  reg [7:0] sc2mac_wt_data28_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1246" *)
  wire [7:0] sc2mac_wt_data29_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1508" *)
  reg [7:0] sc2mac_wt_data29_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1247" *)
  wire [7:0] sc2mac_wt_data2_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1509" *)
  reg [7:0] sc2mac_wt_data2_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1248" *)
  wire [7:0] sc2mac_wt_data30_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1510" *)
  reg [7:0] sc2mac_wt_data30_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1249" *)
  wire [7:0] sc2mac_wt_data31_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1511" *)
  reg [7:0] sc2mac_wt_data31_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1250" *)
  wire [7:0] sc2mac_wt_data32_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1512" *)
  reg [7:0] sc2mac_wt_data32_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1251" *)
  wire [7:0] sc2mac_wt_data33_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1513" *)
  reg [7:0] sc2mac_wt_data33_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1252" *)
  wire [7:0] sc2mac_wt_data34_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1514" *)
  reg [7:0] sc2mac_wt_data34_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1253" *)
  wire [7:0] sc2mac_wt_data35_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1515" *)
  reg [7:0] sc2mac_wt_data35_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1254" *)
  wire [7:0] sc2mac_wt_data36_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1516" *)
  reg [7:0] sc2mac_wt_data36_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1255" *)
  wire [7:0] sc2mac_wt_data37_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1517" *)
  reg [7:0] sc2mac_wt_data37_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1256" *)
  wire [7:0] sc2mac_wt_data38_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1518" *)
  reg [7:0] sc2mac_wt_data38_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1257" *)
  wire [7:0] sc2mac_wt_data39_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1519" *)
  reg [7:0] sc2mac_wt_data39_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1258" *)
  wire [7:0] sc2mac_wt_data3_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1520" *)
  reg [7:0] sc2mac_wt_data3_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1259" *)
  wire [7:0] sc2mac_wt_data40_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1521" *)
  reg [7:0] sc2mac_wt_data40_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1260" *)
  wire [7:0] sc2mac_wt_data41_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1522" *)
  reg [7:0] sc2mac_wt_data41_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1261" *)
  wire [7:0] sc2mac_wt_data42_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1523" *)
  reg [7:0] sc2mac_wt_data42_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1262" *)
  wire [7:0] sc2mac_wt_data43_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1524" *)
  reg [7:0] sc2mac_wt_data43_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1263" *)
  wire [7:0] sc2mac_wt_data44_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1525" *)
  reg [7:0] sc2mac_wt_data44_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1264" *)
  wire [7:0] sc2mac_wt_data45_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1526" *)
  reg [7:0] sc2mac_wt_data45_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1265" *)
  wire [7:0] sc2mac_wt_data46_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1527" *)
  reg [7:0] sc2mac_wt_data46_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1266" *)
  wire [7:0] sc2mac_wt_data47_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1528" *)
  reg [7:0] sc2mac_wt_data47_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1267" *)
  wire [7:0] sc2mac_wt_data48_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1529" *)
  reg [7:0] sc2mac_wt_data48_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1268" *)
  wire [7:0] sc2mac_wt_data49_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1530" *)
  reg [7:0] sc2mac_wt_data49_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1269" *)
  wire [7:0] sc2mac_wt_data4_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1531" *)
  reg [7:0] sc2mac_wt_data4_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1270" *)
  wire [7:0] sc2mac_wt_data50_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1532" *)
  reg [7:0] sc2mac_wt_data50_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1271" *)
  wire [7:0] sc2mac_wt_data51_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1533" *)
  reg [7:0] sc2mac_wt_data51_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1272" *)
  wire [7:0] sc2mac_wt_data52_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1534" *)
  reg [7:0] sc2mac_wt_data52_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1273" *)
  wire [7:0] sc2mac_wt_data53_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1535" *)
  reg [7:0] sc2mac_wt_data53_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1274" *)
  wire [7:0] sc2mac_wt_data54_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1536" *)
  reg [7:0] sc2mac_wt_data54_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1275" *)
  wire [7:0] sc2mac_wt_data55_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1537" *)
  reg [7:0] sc2mac_wt_data55_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1276" *)
  wire [7:0] sc2mac_wt_data56_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1538" *)
  reg [7:0] sc2mac_wt_data56_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1277" *)
  wire [7:0] sc2mac_wt_data57_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1539" *)
  reg [7:0] sc2mac_wt_data57_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1278" *)
  wire [7:0] sc2mac_wt_data58_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1540" *)
  reg [7:0] sc2mac_wt_data58_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1279" *)
  wire [7:0] sc2mac_wt_data59_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1541" *)
  reg [7:0] sc2mac_wt_data59_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1280" *)
  wire [7:0] sc2mac_wt_data5_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1542" *)
  reg [7:0] sc2mac_wt_data5_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1281" *)
  wire [7:0] sc2mac_wt_data60_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1543" *)
  reg [7:0] sc2mac_wt_data60_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1282" *)
  wire [7:0] sc2mac_wt_data61_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1544" *)
  reg [7:0] sc2mac_wt_data61_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1283" *)
  wire [7:0] sc2mac_wt_data62_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1545" *)
  reg [7:0] sc2mac_wt_data62_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1284" *)
  wire [7:0] sc2mac_wt_data63_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1546" *)
  reg [7:0] sc2mac_wt_data63_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1285" *)
  wire [7:0] sc2mac_wt_data64_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1547" *)
  reg [7:0] sc2mac_wt_data64_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1286" *)
  wire [7:0] sc2mac_wt_data65_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1548" *)
  reg [7:0] sc2mac_wt_data65_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1287" *)
  wire [7:0] sc2mac_wt_data66_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1549" *)
  reg [7:0] sc2mac_wt_data66_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1288" *)
  wire [7:0] sc2mac_wt_data67_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1550" *)
  reg [7:0] sc2mac_wt_data67_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1289" *)
  wire [7:0] sc2mac_wt_data68_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1551" *)
  reg [7:0] sc2mac_wt_data68_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1290" *)
  wire [7:0] sc2mac_wt_data69_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1552" *)
  reg [7:0] sc2mac_wt_data69_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1291" *)
  wire [7:0] sc2mac_wt_data6_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1553" *)
  reg [7:0] sc2mac_wt_data6_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1292" *)
  wire [7:0] sc2mac_wt_data70_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1554" *)
  reg [7:0] sc2mac_wt_data70_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1293" *)
  wire [7:0] sc2mac_wt_data71_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1555" *)
  reg [7:0] sc2mac_wt_data71_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1294" *)
  wire [7:0] sc2mac_wt_data72_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1556" *)
  reg [7:0] sc2mac_wt_data72_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1295" *)
  wire [7:0] sc2mac_wt_data73_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1557" *)
  reg [7:0] sc2mac_wt_data73_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1296" *)
  wire [7:0] sc2mac_wt_data74_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1558" *)
  reg [7:0] sc2mac_wt_data74_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1297" *)
  wire [7:0] sc2mac_wt_data75_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1559" *)
  reg [7:0] sc2mac_wt_data75_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1298" *)
  wire [7:0] sc2mac_wt_data76_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1560" *)
  reg [7:0] sc2mac_wt_data76_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1299" *)
  wire [7:0] sc2mac_wt_data77_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1561" *)
  reg [7:0] sc2mac_wt_data77_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1300" *)
  wire [7:0] sc2mac_wt_data78_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1562" *)
  reg [7:0] sc2mac_wt_data78_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1301" *)
  wire [7:0] sc2mac_wt_data79_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1563" *)
  reg [7:0] sc2mac_wt_data79_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1302" *)
  wire [7:0] sc2mac_wt_data7_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1564" *)
  reg [7:0] sc2mac_wt_data7_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1303" *)
  wire [7:0] sc2mac_wt_data80_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1565" *)
  reg [7:0] sc2mac_wt_data80_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1304" *)
  wire [7:0] sc2mac_wt_data81_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1566" *)
  reg [7:0] sc2mac_wt_data81_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1305" *)
  wire [7:0] sc2mac_wt_data82_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1567" *)
  reg [7:0] sc2mac_wt_data82_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1306" *)
  wire [7:0] sc2mac_wt_data83_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1568" *)
  reg [7:0] sc2mac_wt_data83_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1307" *)
  wire [7:0] sc2mac_wt_data84_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1569" *)
  reg [7:0] sc2mac_wt_data84_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1308" *)
  wire [7:0] sc2mac_wt_data85_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1570" *)
  reg [7:0] sc2mac_wt_data85_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1309" *)
  wire [7:0] sc2mac_wt_data86_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1571" *)
  reg [7:0] sc2mac_wt_data86_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1310" *)
  wire [7:0] sc2mac_wt_data87_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1572" *)
  reg [7:0] sc2mac_wt_data87_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1311" *)
  wire [7:0] sc2mac_wt_data88_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1573" *)
  reg [7:0] sc2mac_wt_data88_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1312" *)
  wire [7:0] sc2mac_wt_data89_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1574" *)
  reg [7:0] sc2mac_wt_data89_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1313" *)
  wire [7:0] sc2mac_wt_data8_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1575" *)
  reg [7:0] sc2mac_wt_data8_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1314" *)
  wire [7:0] sc2mac_wt_data90_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1576" *)
  reg [7:0] sc2mac_wt_data90_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1315" *)
  wire [7:0] sc2mac_wt_data91_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1577" *)
  reg [7:0] sc2mac_wt_data91_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1316" *)
  wire [7:0] sc2mac_wt_data92_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1578" *)
  reg [7:0] sc2mac_wt_data92_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1317" *)
  wire [7:0] sc2mac_wt_data93_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1579" *)
  reg [7:0] sc2mac_wt_data93_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1318" *)
  wire [7:0] sc2mac_wt_data94_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1580" *)
  reg [7:0] sc2mac_wt_data94_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1319" *)
  wire [7:0] sc2mac_wt_data95_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1581" *)
  reg [7:0] sc2mac_wt_data95_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1320" *)
  wire [7:0] sc2mac_wt_data96_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1582" *)
  reg [7:0] sc2mac_wt_data96_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1321" *)
  wire [7:0] sc2mac_wt_data97_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1583" *)
  reg [7:0] sc2mac_wt_data97_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1322" *)
  wire [7:0] sc2mac_wt_data98_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1584" *)
  reg [7:0] sc2mac_wt_data98_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1323" *)
  wire [7:0] sc2mac_wt_data99_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1585" *)
  reg [7:0] sc2mac_wt_data99_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1324" *)
  wire [7:0] sc2mac_wt_data9_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1586" *)
  reg [7:0] sc2mac_wt_data9_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:806" *)
  output [7:0] sc2mac_wt_dst_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:807" *)
  output [7:0] sc2mac_wt_dst_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:816" *)
  output [7:0] sc2mac_wt_dst_data10;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:906" *)
  output [7:0] sc2mac_wt_dst_data100;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:907" *)
  output [7:0] sc2mac_wt_dst_data101;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:908" *)
  output [7:0] sc2mac_wt_dst_data102;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:909" *)
  output [7:0] sc2mac_wt_dst_data103;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:910" *)
  output [7:0] sc2mac_wt_dst_data104;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:911" *)
  output [7:0] sc2mac_wt_dst_data105;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:912" *)
  output [7:0] sc2mac_wt_dst_data106;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:913" *)
  output [7:0] sc2mac_wt_dst_data107;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:914" *)
  output [7:0] sc2mac_wt_dst_data108;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:915" *)
  output [7:0] sc2mac_wt_dst_data109;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:817" *)
  output [7:0] sc2mac_wt_dst_data11;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:916" *)
  output [7:0] sc2mac_wt_dst_data110;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:917" *)
  output [7:0] sc2mac_wt_dst_data111;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:918" *)
  output [7:0] sc2mac_wt_dst_data112;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:919" *)
  output [7:0] sc2mac_wt_dst_data113;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:920" *)
  output [7:0] sc2mac_wt_dst_data114;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:921" *)
  output [7:0] sc2mac_wt_dst_data115;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:922" *)
  output [7:0] sc2mac_wt_dst_data116;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:923" *)
  output [7:0] sc2mac_wt_dst_data117;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:924" *)
  output [7:0] sc2mac_wt_dst_data118;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:925" *)
  output [7:0] sc2mac_wt_dst_data119;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:818" *)
  output [7:0] sc2mac_wt_dst_data12;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:926" *)
  output [7:0] sc2mac_wt_dst_data120;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:927" *)
  output [7:0] sc2mac_wt_dst_data121;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:928" *)
  output [7:0] sc2mac_wt_dst_data122;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:929" *)
  output [7:0] sc2mac_wt_dst_data123;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:930" *)
  output [7:0] sc2mac_wt_dst_data124;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:931" *)
  output [7:0] sc2mac_wt_dst_data125;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:932" *)
  output [7:0] sc2mac_wt_dst_data126;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:933" *)
  output [7:0] sc2mac_wt_dst_data127;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:819" *)
  output [7:0] sc2mac_wt_dst_data13;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:820" *)
  output [7:0] sc2mac_wt_dst_data14;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:821" *)
  output [7:0] sc2mac_wt_dst_data15;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:822" *)
  output [7:0] sc2mac_wt_dst_data16;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:823" *)
  output [7:0] sc2mac_wt_dst_data17;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:824" *)
  output [7:0] sc2mac_wt_dst_data18;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:825" *)
  output [7:0] sc2mac_wt_dst_data19;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:808" *)
  output [7:0] sc2mac_wt_dst_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:826" *)
  output [7:0] sc2mac_wt_dst_data20;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:827" *)
  output [7:0] sc2mac_wt_dst_data21;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:828" *)
  output [7:0] sc2mac_wt_dst_data22;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:829" *)
  output [7:0] sc2mac_wt_dst_data23;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:830" *)
  output [7:0] sc2mac_wt_dst_data24;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:831" *)
  output [7:0] sc2mac_wt_dst_data25;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:832" *)
  output [7:0] sc2mac_wt_dst_data26;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:833" *)
  output [7:0] sc2mac_wt_dst_data27;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:834" *)
  output [7:0] sc2mac_wt_dst_data28;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:835" *)
  output [7:0] sc2mac_wt_dst_data29;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:809" *)
  output [7:0] sc2mac_wt_dst_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:836" *)
  output [7:0] sc2mac_wt_dst_data30;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:837" *)
  output [7:0] sc2mac_wt_dst_data31;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:838" *)
  output [7:0] sc2mac_wt_dst_data32;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:839" *)
  output [7:0] sc2mac_wt_dst_data33;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:840" *)
  output [7:0] sc2mac_wt_dst_data34;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:841" *)
  output [7:0] sc2mac_wt_dst_data35;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:842" *)
  output [7:0] sc2mac_wt_dst_data36;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:843" *)
  output [7:0] sc2mac_wt_dst_data37;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:844" *)
  output [7:0] sc2mac_wt_dst_data38;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:845" *)
  output [7:0] sc2mac_wt_dst_data39;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:810" *)
  output [7:0] sc2mac_wt_dst_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:846" *)
  output [7:0] sc2mac_wt_dst_data40;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:847" *)
  output [7:0] sc2mac_wt_dst_data41;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:848" *)
  output [7:0] sc2mac_wt_dst_data42;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:849" *)
  output [7:0] sc2mac_wt_dst_data43;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:850" *)
  output [7:0] sc2mac_wt_dst_data44;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:851" *)
  output [7:0] sc2mac_wt_dst_data45;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:852" *)
  output [7:0] sc2mac_wt_dst_data46;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:853" *)
  output [7:0] sc2mac_wt_dst_data47;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:854" *)
  output [7:0] sc2mac_wt_dst_data48;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:855" *)
  output [7:0] sc2mac_wt_dst_data49;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:811" *)
  output [7:0] sc2mac_wt_dst_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:856" *)
  output [7:0] sc2mac_wt_dst_data50;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:857" *)
  output [7:0] sc2mac_wt_dst_data51;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:858" *)
  output [7:0] sc2mac_wt_dst_data52;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:859" *)
  output [7:0] sc2mac_wt_dst_data53;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:860" *)
  output [7:0] sc2mac_wt_dst_data54;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:861" *)
  output [7:0] sc2mac_wt_dst_data55;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:862" *)
  output [7:0] sc2mac_wt_dst_data56;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:863" *)
  output [7:0] sc2mac_wt_dst_data57;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:864" *)
  output [7:0] sc2mac_wt_dst_data58;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:865" *)
  output [7:0] sc2mac_wt_dst_data59;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:812" *)
  output [7:0] sc2mac_wt_dst_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:866" *)
  output [7:0] sc2mac_wt_dst_data60;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:867" *)
  output [7:0] sc2mac_wt_dst_data61;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:868" *)
  output [7:0] sc2mac_wt_dst_data62;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:869" *)
  output [7:0] sc2mac_wt_dst_data63;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:870" *)
  output [7:0] sc2mac_wt_dst_data64;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:871" *)
  output [7:0] sc2mac_wt_dst_data65;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:872" *)
  output [7:0] sc2mac_wt_dst_data66;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:873" *)
  output [7:0] sc2mac_wt_dst_data67;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:874" *)
  output [7:0] sc2mac_wt_dst_data68;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:875" *)
  output [7:0] sc2mac_wt_dst_data69;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:813" *)
  output [7:0] sc2mac_wt_dst_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:876" *)
  output [7:0] sc2mac_wt_dst_data70;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:877" *)
  output [7:0] sc2mac_wt_dst_data71;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:878" *)
  output [7:0] sc2mac_wt_dst_data72;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:879" *)
  output [7:0] sc2mac_wt_dst_data73;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:880" *)
  output [7:0] sc2mac_wt_dst_data74;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:881" *)
  output [7:0] sc2mac_wt_dst_data75;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:882" *)
  output [7:0] sc2mac_wt_dst_data76;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:883" *)
  output [7:0] sc2mac_wt_dst_data77;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:884" *)
  output [7:0] sc2mac_wt_dst_data78;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:885" *)
  output [7:0] sc2mac_wt_dst_data79;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:814" *)
  output [7:0] sc2mac_wt_dst_data8;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:886" *)
  output [7:0] sc2mac_wt_dst_data80;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:887" *)
  output [7:0] sc2mac_wt_dst_data81;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:888" *)
  output [7:0] sc2mac_wt_dst_data82;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:889" *)
  output [7:0] sc2mac_wt_dst_data83;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:890" *)
  output [7:0] sc2mac_wt_dst_data84;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:891" *)
  output [7:0] sc2mac_wt_dst_data85;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:892" *)
  output [7:0] sc2mac_wt_dst_data86;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:893" *)
  output [7:0] sc2mac_wt_dst_data87;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:894" *)
  output [7:0] sc2mac_wt_dst_data88;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:895" *)
  output [7:0] sc2mac_wt_dst_data89;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:815" *)
  output [7:0] sc2mac_wt_dst_data9;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:896" *)
  output [7:0] sc2mac_wt_dst_data90;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:897" *)
  output [7:0] sc2mac_wt_dst_data91;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:898" *)
  output [7:0] sc2mac_wt_dst_data92;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:899" *)
  output [7:0] sc2mac_wt_dst_data93;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:900" *)
  output [7:0] sc2mac_wt_dst_data94;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:901" *)
  output [7:0] sc2mac_wt_dst_data95;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:902" *)
  output [7:0] sc2mac_wt_dst_data96;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:903" *)
  output [7:0] sc2mac_wt_dst_data97;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:904" *)
  output [7:0] sc2mac_wt_dst_data98;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:905" *)
  output [7:0] sc2mac_wt_dst_data99;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:805" *)
  output [127:0] sc2mac_wt_dst_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:804" *)
  output sc2mac_wt_dst_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:934" *)
  output [7:0] sc2mac_wt_dst_sel;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1325" *)
  wire [127:0] sc2mac_wt_mask_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1587" *)
  reg [127:0] sc2mac_wt_mask_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1326" *)
  wire sc2mac_wt_pvld_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1588" *)
  reg sc2mac_wt_pvld_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1327" *)
  wire [7:0] sc2mac_wt_sel_d0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1589" *)
  reg [7:0] sc2mac_wt_sel_d1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:544" *)
  input [7:0] sc2mac_wt_src_data0;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:545" *)
  input [7:0] sc2mac_wt_src_data1;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:554" *)
  input [7:0] sc2mac_wt_src_data10;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:644" *)
  input [7:0] sc2mac_wt_src_data100;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:645" *)
  input [7:0] sc2mac_wt_src_data101;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:646" *)
  input [7:0] sc2mac_wt_src_data102;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:647" *)
  input [7:0] sc2mac_wt_src_data103;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:648" *)
  input [7:0] sc2mac_wt_src_data104;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:649" *)
  input [7:0] sc2mac_wt_src_data105;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:650" *)
  input [7:0] sc2mac_wt_src_data106;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:651" *)
  input [7:0] sc2mac_wt_src_data107;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:652" *)
  input [7:0] sc2mac_wt_src_data108;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:653" *)
  input [7:0] sc2mac_wt_src_data109;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:555" *)
  input [7:0] sc2mac_wt_src_data11;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:654" *)
  input [7:0] sc2mac_wt_src_data110;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:655" *)
  input [7:0] sc2mac_wt_src_data111;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:656" *)
  input [7:0] sc2mac_wt_src_data112;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:657" *)
  input [7:0] sc2mac_wt_src_data113;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:658" *)
  input [7:0] sc2mac_wt_src_data114;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:659" *)
  input [7:0] sc2mac_wt_src_data115;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:660" *)
  input [7:0] sc2mac_wt_src_data116;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:661" *)
  input [7:0] sc2mac_wt_src_data117;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:662" *)
  input [7:0] sc2mac_wt_src_data118;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:663" *)
  input [7:0] sc2mac_wt_src_data119;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:556" *)
  input [7:0] sc2mac_wt_src_data12;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:664" *)
  input [7:0] sc2mac_wt_src_data120;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:665" *)
  input [7:0] sc2mac_wt_src_data121;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:666" *)
  input [7:0] sc2mac_wt_src_data122;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:667" *)
  input [7:0] sc2mac_wt_src_data123;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:668" *)
  input [7:0] sc2mac_wt_src_data124;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:669" *)
  input [7:0] sc2mac_wt_src_data125;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:670" *)
  input [7:0] sc2mac_wt_src_data126;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:671" *)
  input [7:0] sc2mac_wt_src_data127;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:557" *)
  input [7:0] sc2mac_wt_src_data13;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:558" *)
  input [7:0] sc2mac_wt_src_data14;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:559" *)
  input [7:0] sc2mac_wt_src_data15;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:560" *)
  input [7:0] sc2mac_wt_src_data16;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:561" *)
  input [7:0] sc2mac_wt_src_data17;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:562" *)
  input [7:0] sc2mac_wt_src_data18;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:563" *)
  input [7:0] sc2mac_wt_src_data19;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:546" *)
  input [7:0] sc2mac_wt_src_data2;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:564" *)
  input [7:0] sc2mac_wt_src_data20;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:565" *)
  input [7:0] sc2mac_wt_src_data21;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:566" *)
  input [7:0] sc2mac_wt_src_data22;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:567" *)
  input [7:0] sc2mac_wt_src_data23;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:568" *)
  input [7:0] sc2mac_wt_src_data24;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:569" *)
  input [7:0] sc2mac_wt_src_data25;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:570" *)
  input [7:0] sc2mac_wt_src_data26;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:571" *)
  input [7:0] sc2mac_wt_src_data27;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:572" *)
  input [7:0] sc2mac_wt_src_data28;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:573" *)
  input [7:0] sc2mac_wt_src_data29;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:547" *)
  input [7:0] sc2mac_wt_src_data3;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:574" *)
  input [7:0] sc2mac_wt_src_data30;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:575" *)
  input [7:0] sc2mac_wt_src_data31;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:576" *)
  input [7:0] sc2mac_wt_src_data32;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:577" *)
  input [7:0] sc2mac_wt_src_data33;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:578" *)
  input [7:0] sc2mac_wt_src_data34;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:579" *)
  input [7:0] sc2mac_wt_src_data35;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:580" *)
  input [7:0] sc2mac_wt_src_data36;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:581" *)
  input [7:0] sc2mac_wt_src_data37;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:582" *)
  input [7:0] sc2mac_wt_src_data38;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:583" *)
  input [7:0] sc2mac_wt_src_data39;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:548" *)
  input [7:0] sc2mac_wt_src_data4;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:584" *)
  input [7:0] sc2mac_wt_src_data40;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:585" *)
  input [7:0] sc2mac_wt_src_data41;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:586" *)
  input [7:0] sc2mac_wt_src_data42;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:587" *)
  input [7:0] sc2mac_wt_src_data43;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:588" *)
  input [7:0] sc2mac_wt_src_data44;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:589" *)
  input [7:0] sc2mac_wt_src_data45;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:590" *)
  input [7:0] sc2mac_wt_src_data46;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:591" *)
  input [7:0] sc2mac_wt_src_data47;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:592" *)
  input [7:0] sc2mac_wt_src_data48;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:593" *)
  input [7:0] sc2mac_wt_src_data49;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:549" *)
  input [7:0] sc2mac_wt_src_data5;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:594" *)
  input [7:0] sc2mac_wt_src_data50;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:595" *)
  input [7:0] sc2mac_wt_src_data51;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:596" *)
  input [7:0] sc2mac_wt_src_data52;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:597" *)
  input [7:0] sc2mac_wt_src_data53;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:598" *)
  input [7:0] sc2mac_wt_src_data54;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:599" *)
  input [7:0] sc2mac_wt_src_data55;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:600" *)
  input [7:0] sc2mac_wt_src_data56;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:601" *)
  input [7:0] sc2mac_wt_src_data57;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:602" *)
  input [7:0] sc2mac_wt_src_data58;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:603" *)
  input [7:0] sc2mac_wt_src_data59;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:550" *)
  input [7:0] sc2mac_wt_src_data6;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:604" *)
  input [7:0] sc2mac_wt_src_data60;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:605" *)
  input [7:0] sc2mac_wt_src_data61;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:606" *)
  input [7:0] sc2mac_wt_src_data62;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:607" *)
  input [7:0] sc2mac_wt_src_data63;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:608" *)
  input [7:0] sc2mac_wt_src_data64;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:609" *)
  input [7:0] sc2mac_wt_src_data65;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:610" *)
  input [7:0] sc2mac_wt_src_data66;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:611" *)
  input [7:0] sc2mac_wt_src_data67;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:612" *)
  input [7:0] sc2mac_wt_src_data68;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:613" *)
  input [7:0] sc2mac_wt_src_data69;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:551" *)
  input [7:0] sc2mac_wt_src_data7;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:614" *)
  input [7:0] sc2mac_wt_src_data70;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:615" *)
  input [7:0] sc2mac_wt_src_data71;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:616" *)
  input [7:0] sc2mac_wt_src_data72;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:617" *)
  input [7:0] sc2mac_wt_src_data73;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:618" *)
  input [7:0] sc2mac_wt_src_data74;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:619" *)
  input [7:0] sc2mac_wt_src_data75;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:620" *)
  input [7:0] sc2mac_wt_src_data76;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:621" *)
  input [7:0] sc2mac_wt_src_data77;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:622" *)
  input [7:0] sc2mac_wt_src_data78;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:623" *)
  input [7:0] sc2mac_wt_src_data79;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:552" *)
  input [7:0] sc2mac_wt_src_data8;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:624" *)
  input [7:0] sc2mac_wt_src_data80;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:625" *)
  input [7:0] sc2mac_wt_src_data81;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:626" *)
  input [7:0] sc2mac_wt_src_data82;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:627" *)
  input [7:0] sc2mac_wt_src_data83;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:628" *)
  input [7:0] sc2mac_wt_src_data84;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:629" *)
  input [7:0] sc2mac_wt_src_data85;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:630" *)
  input [7:0] sc2mac_wt_src_data86;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:631" *)
  input [7:0] sc2mac_wt_src_data87;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:632" *)
  input [7:0] sc2mac_wt_src_data88;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:633" *)
  input [7:0] sc2mac_wt_src_data89;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:553" *)
  input [7:0] sc2mac_wt_src_data9;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:634" *)
  input [7:0] sc2mac_wt_src_data90;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:635" *)
  input [7:0] sc2mac_wt_src_data91;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:636" *)
  input [7:0] sc2mac_wt_src_data92;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:637" *)
  input [7:0] sc2mac_wt_src_data93;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:638" *)
  input [7:0] sc2mac_wt_src_data94;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:639" *)
  input [7:0] sc2mac_wt_src_data95;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:640" *)
  input [7:0] sc2mac_wt_src_data96;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:641" *)
  input [7:0] sc2mac_wt_src_data97;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:642" *)
  input [7:0] sc2mac_wt_src_data98;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:643" *)
  input [7:0] sc2mac_wt_src_data99;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:543" *)
  input [127:0] sc2mac_wt_src_mask;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:542" *)
  input sc2mac_wt_src_pvld;
  (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:672" *)
  input [7:0] sc2mac_wt_src_sel;
  assign _260_ = sc2mac_wt_src_pvld | (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1863" *) sc2mac_wt_pvld_d1;
  assign _261_ = sc2mac_dat_src_pvld | (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3272" *) sc2mac_dat_pvld_d1;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data127_d1 <= _030_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data126_d1 <= _029_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data125_d1 <= _028_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data124_d1 <= _027_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data123_d1 <= _026_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data122_d1 <= _025_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data121_d1 <= _024_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data120_d1 <= _023_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data119_d1 <= _021_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data118_d1 <= _020_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data117_d1 <= _019_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data116_d1 <= _018_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data115_d1 <= _017_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data114_d1 <= _016_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data113_d1 <= _015_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data112_d1 <= _014_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data111_d1 <= _013_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data110_d1 <= _012_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data109_d1 <= _010_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data108_d1 <= _009_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data107_d1 <= _008_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data106_d1 <= _007_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data105_d1 <= _006_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data104_d1 <= _005_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data103_d1 <= _004_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data102_d1 <= _003_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data101_d1 <= _002_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data100_d1 <= _001_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data99_d1 <= _126_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data98_d1 <= _125_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data97_d1 <= _124_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data96_d1 <= _123_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data95_d1 <= _122_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data94_d1 <= _121_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data93_d1 <= _120_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data92_d1 <= _119_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data91_d1 <= _118_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data90_d1 <= _117_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data89_d1 <= _115_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data88_d1 <= _114_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data87_d1 <= _113_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data86_d1 <= _112_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data85_d1 <= _111_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data84_d1 <= _110_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data83_d1 <= _109_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data82_d1 <= _108_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data81_d1 <= _107_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data80_d1 <= _106_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data79_d1 <= _104_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data78_d1 <= _103_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data77_d1 <= _102_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data76_d1 <= _101_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data75_d1 <= _100_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data74_d1 <= _099_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data73_d1 <= _098_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data72_d1 <= _097_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data71_d1 <= _096_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data70_d1 <= _095_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data69_d1 <= _093_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data68_d1 <= _092_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data67_d1 <= _091_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data66_d1 <= _090_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data65_d1 <= _089_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data64_d1 <= _088_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data63_d1 <= _087_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data62_d1 <= _086_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data61_d1 <= _085_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data60_d1 <= _084_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data59_d1 <= _082_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data58_d1 <= _081_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data57_d1 <= _080_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data56_d1 <= _079_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data55_d1 <= _078_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data54_d1 <= _077_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data53_d1 <= _076_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data52_d1 <= _075_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data51_d1 <= _074_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data50_d1 <= _073_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data49_d1 <= _071_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data48_d1 <= _070_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data47_d1 <= _069_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data46_d1 <= _068_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data45_d1 <= _067_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data44_d1 <= _066_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data43_d1 <= _065_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data42_d1 <= _064_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data41_d1 <= _063_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data40_d1 <= _062_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data39_d1 <= _060_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data38_d1 <= _059_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data37_d1 <= _058_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data36_d1 <= _057_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data35_d1 <= _056_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data34_d1 <= _055_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data33_d1 <= _054_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data32_d1 <= _053_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data31_d1 <= _052_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data30_d1 <= _051_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data29_d1 <= _049_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data28_d1 <= _048_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data27_d1 <= _047_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data26_d1 <= _046_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data25_d1 <= _045_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data24_d1 <= _044_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data23_d1 <= _043_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data22_d1 <= _042_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data21_d1 <= _041_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data20_d1 <= _040_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data19_d1 <= _038_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data18_d1 <= _037_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data17_d1 <= _036_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data16_d1 <= _035_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data15_d1 <= _034_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data14_d1 <= _033_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data13_d1 <= _032_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data12_d1 <= _031_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data11_d1 <= _022_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data10_d1 <= _011_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data9_d1 <= _127_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data8_d1 <= _116_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data7_d1 <= _105_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data6_d1 <= _094_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data5_d1 <= _083_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data4_d1 <= _072_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data3_d1 <= _061_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data2_d1 <= _050_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data1_d1 <= _039_;
  always @(posedge nvdla_core_clk)
      sc2mac_dat_data0_d1 <= _000_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_mask_d1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      sc2mac_dat_mask_d1 <= _128_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_pd_d1 <= 9'b000000000;
    else
      sc2mac_dat_pd_d1 <= _129_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_dat_pvld_d1 <= 1'b0;
    else
      sc2mac_dat_pvld_d1 <= sc2mac_dat_src_pvld;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data127_d1 <= _160_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data126_d1 <= _159_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data125_d1 <= _158_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data124_d1 <= _157_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data123_d1 <= _156_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data122_d1 <= _155_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data121_d1 <= _154_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data120_d1 <= _153_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data119_d1 <= _151_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data118_d1 <= _150_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data117_d1 <= _149_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data116_d1 <= _148_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data115_d1 <= _147_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data114_d1 <= _146_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data113_d1 <= _145_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data112_d1 <= _144_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data111_d1 <= _143_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data110_d1 <= _142_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data109_d1 <= _140_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data108_d1 <= _139_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data107_d1 <= _138_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data106_d1 <= _137_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data105_d1 <= _136_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data104_d1 <= _135_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data103_d1 <= _134_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data102_d1 <= _133_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data101_d1 <= _132_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data100_d1 <= _131_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data99_d1 <= _256_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data98_d1 <= _255_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data97_d1 <= _254_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data96_d1 <= _253_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data95_d1 <= _252_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data94_d1 <= _251_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data93_d1 <= _250_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data92_d1 <= _249_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data91_d1 <= _248_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data90_d1 <= _247_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data89_d1 <= _245_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data88_d1 <= _244_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data87_d1 <= _243_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data86_d1 <= _242_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data85_d1 <= _241_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data84_d1 <= _240_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data83_d1 <= _239_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data82_d1 <= _238_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data81_d1 <= _237_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data80_d1 <= _236_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data79_d1 <= _234_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data78_d1 <= _233_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data77_d1 <= _232_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data76_d1 <= _231_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data75_d1 <= _230_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data74_d1 <= _229_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data73_d1 <= _228_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data72_d1 <= _227_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data71_d1 <= _226_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data70_d1 <= _225_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data69_d1 <= _223_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data68_d1 <= _222_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data67_d1 <= _221_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data66_d1 <= _220_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data65_d1 <= _219_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data64_d1 <= _218_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data63_d1 <= _217_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data62_d1 <= _216_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data61_d1 <= _215_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data60_d1 <= _214_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data59_d1 <= _212_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data58_d1 <= _211_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data57_d1 <= _210_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data56_d1 <= _209_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data55_d1 <= _208_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data54_d1 <= _207_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data53_d1 <= _206_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data52_d1 <= _205_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data51_d1 <= _204_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data50_d1 <= _203_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data49_d1 <= _201_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data48_d1 <= _200_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data47_d1 <= _199_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data46_d1 <= _198_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data45_d1 <= _197_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data44_d1 <= _196_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data43_d1 <= _195_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data42_d1 <= _194_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data41_d1 <= _193_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data40_d1 <= _192_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data39_d1 <= _190_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data38_d1 <= _189_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data37_d1 <= _188_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data36_d1 <= _187_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data35_d1 <= _186_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data34_d1 <= _185_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data33_d1 <= _184_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data32_d1 <= _183_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data31_d1 <= _182_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data30_d1 <= _181_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data29_d1 <= _179_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data28_d1 <= _178_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data27_d1 <= _177_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data26_d1 <= _176_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data25_d1 <= _175_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data24_d1 <= _174_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data23_d1 <= _173_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data22_d1 <= _172_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data21_d1 <= _171_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data20_d1 <= _170_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data19_d1 <= _168_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data18_d1 <= _167_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data17_d1 <= _166_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data16_d1 <= _165_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data15_d1 <= _164_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data14_d1 <= _163_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data13_d1 <= _162_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data12_d1 <= _161_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data11_d1 <= _152_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data10_d1 <= _141_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data9_d1 <= _257_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data8_d1 <= _246_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data7_d1 <= _235_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data6_d1 <= _224_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data5_d1 <= _213_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data4_d1 <= _202_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data3_d1 <= _191_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data2_d1 <= _180_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data1_d1 <= _169_;
  always @(posedge nvdla_core_clk)
      sc2mac_wt_data0_d1 <= _130_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_wt_mask_d1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      sc2mac_wt_mask_d1 <= _258_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_wt_sel_d1 <= 8'b00000000;
    else
      sc2mac_wt_sel_d1 <= _259_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sc2mac_wt_pvld_d1 <= 1'b0;
    else
      sc2mac_wt_pvld_d1 <= sc2mac_wt_src_pvld;
  assign _030_ = sc2mac_dat_src_mask[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4661" *) sc2mac_dat_src_data127 : sc2mac_dat_data127_d1;
  assign _029_ = sc2mac_dat_src_mask[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4651" *) sc2mac_dat_src_data126 : sc2mac_dat_data126_d1;
  assign _028_ = sc2mac_dat_src_mask[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4641" *) sc2mac_dat_src_data125 : sc2mac_dat_data125_d1;
  assign _027_ = sc2mac_dat_src_mask[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4631" *) sc2mac_dat_src_data124 : sc2mac_dat_data124_d1;
  assign _026_ = sc2mac_dat_src_mask[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4621" *) sc2mac_dat_src_data123 : sc2mac_dat_data123_d1;
  assign _025_ = sc2mac_dat_src_mask[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4611" *) sc2mac_dat_src_data122 : sc2mac_dat_data122_d1;
  assign _024_ = sc2mac_dat_src_mask[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4601" *) sc2mac_dat_src_data121 : sc2mac_dat_data121_d1;
  assign _023_ = sc2mac_dat_src_mask[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4591" *) sc2mac_dat_src_data120 : sc2mac_dat_data120_d1;
  assign _021_ = sc2mac_dat_src_mask[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4581" *) sc2mac_dat_src_data119 : sc2mac_dat_data119_d1;
  assign _020_ = sc2mac_dat_src_mask[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4571" *) sc2mac_dat_src_data118 : sc2mac_dat_data118_d1;
  assign _019_ = sc2mac_dat_src_mask[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4561" *) sc2mac_dat_src_data117 : sc2mac_dat_data117_d1;
  assign _018_ = sc2mac_dat_src_mask[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4551" *) sc2mac_dat_src_data116 : sc2mac_dat_data116_d1;
  assign _017_ = sc2mac_dat_src_mask[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4541" *) sc2mac_dat_src_data115 : sc2mac_dat_data115_d1;
  assign _016_ = sc2mac_dat_src_mask[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4531" *) sc2mac_dat_src_data114 : sc2mac_dat_data114_d1;
  assign _015_ = sc2mac_dat_src_mask[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4521" *) sc2mac_dat_src_data113 : sc2mac_dat_data113_d1;
  assign _014_ = sc2mac_dat_src_mask[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4511" *) sc2mac_dat_src_data112 : sc2mac_dat_data112_d1;
  assign _013_ = sc2mac_dat_src_mask[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4501" *) sc2mac_dat_src_data111 : sc2mac_dat_data111_d1;
  assign _012_ = sc2mac_dat_src_mask[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4491" *) sc2mac_dat_src_data110 : sc2mac_dat_data110_d1;
  assign _010_ = sc2mac_dat_src_mask[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4481" *) sc2mac_dat_src_data109 : sc2mac_dat_data109_d1;
  assign _009_ = sc2mac_dat_src_mask[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4471" *) sc2mac_dat_src_data108 : sc2mac_dat_data108_d1;
  assign _008_ = sc2mac_dat_src_mask[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4461" *) sc2mac_dat_src_data107 : sc2mac_dat_data107_d1;
  assign _007_ = sc2mac_dat_src_mask[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4451" *) sc2mac_dat_src_data106 : sc2mac_dat_data106_d1;
  assign _006_ = sc2mac_dat_src_mask[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4441" *) sc2mac_dat_src_data105 : sc2mac_dat_data105_d1;
  assign _005_ = sc2mac_dat_src_mask[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4431" *) sc2mac_dat_src_data104 : sc2mac_dat_data104_d1;
  assign _004_ = sc2mac_dat_src_mask[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4421" *) sc2mac_dat_src_data103 : sc2mac_dat_data103_d1;
  assign _003_ = sc2mac_dat_src_mask[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4411" *) sc2mac_dat_src_data102 : sc2mac_dat_data102_d1;
  assign _002_ = sc2mac_dat_src_mask[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4401" *) sc2mac_dat_src_data101 : sc2mac_dat_data101_d1;
  assign _001_ = sc2mac_dat_src_mask[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4391" *) sc2mac_dat_src_data100 : sc2mac_dat_data100_d1;
  assign _126_ = sc2mac_dat_src_mask[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4381" *) sc2mac_dat_src_data99 : sc2mac_dat_data99_d1;
  assign _125_ = sc2mac_dat_src_mask[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4371" *) sc2mac_dat_src_data98 : sc2mac_dat_data98_d1;
  assign _124_ = sc2mac_dat_src_mask[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4361" *) sc2mac_dat_src_data97 : sc2mac_dat_data97_d1;
  assign _123_ = sc2mac_dat_src_mask[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4351" *) sc2mac_dat_src_data96 : sc2mac_dat_data96_d1;
  assign _122_ = sc2mac_dat_src_mask[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4341" *) sc2mac_dat_src_data95 : sc2mac_dat_data95_d1;
  assign _121_ = sc2mac_dat_src_mask[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4331" *) sc2mac_dat_src_data94 : sc2mac_dat_data94_d1;
  assign _120_ = sc2mac_dat_src_mask[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4321" *) sc2mac_dat_src_data93 : sc2mac_dat_data93_d1;
  assign _119_ = sc2mac_dat_src_mask[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4311" *) sc2mac_dat_src_data92 : sc2mac_dat_data92_d1;
  assign _118_ = sc2mac_dat_src_mask[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4301" *) sc2mac_dat_src_data91 : sc2mac_dat_data91_d1;
  assign _117_ = sc2mac_dat_src_mask[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4291" *) sc2mac_dat_src_data90 : sc2mac_dat_data90_d1;
  assign _115_ = sc2mac_dat_src_mask[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4281" *) sc2mac_dat_src_data89 : sc2mac_dat_data89_d1;
  assign _114_ = sc2mac_dat_src_mask[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4271" *) sc2mac_dat_src_data88 : sc2mac_dat_data88_d1;
  assign _113_ = sc2mac_dat_src_mask[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4261" *) sc2mac_dat_src_data87 : sc2mac_dat_data87_d1;
  assign _112_ = sc2mac_dat_src_mask[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4251" *) sc2mac_dat_src_data86 : sc2mac_dat_data86_d1;
  assign _111_ = sc2mac_dat_src_mask[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4241" *) sc2mac_dat_src_data85 : sc2mac_dat_data85_d1;
  assign _110_ = sc2mac_dat_src_mask[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4231" *) sc2mac_dat_src_data84 : sc2mac_dat_data84_d1;
  assign _109_ = sc2mac_dat_src_mask[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4221" *) sc2mac_dat_src_data83 : sc2mac_dat_data83_d1;
  assign _108_ = sc2mac_dat_src_mask[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4211" *) sc2mac_dat_src_data82 : sc2mac_dat_data82_d1;
  assign _107_ = sc2mac_dat_src_mask[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4201" *) sc2mac_dat_src_data81 : sc2mac_dat_data81_d1;
  assign _106_ = sc2mac_dat_src_mask[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4191" *) sc2mac_dat_src_data80 : sc2mac_dat_data80_d1;
  assign _104_ = sc2mac_dat_src_mask[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4181" *) sc2mac_dat_src_data79 : sc2mac_dat_data79_d1;
  assign _103_ = sc2mac_dat_src_mask[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4171" *) sc2mac_dat_src_data78 : sc2mac_dat_data78_d1;
  assign _102_ = sc2mac_dat_src_mask[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4161" *) sc2mac_dat_src_data77 : sc2mac_dat_data77_d1;
  assign _101_ = sc2mac_dat_src_mask[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4151" *) sc2mac_dat_src_data76 : sc2mac_dat_data76_d1;
  assign _100_ = sc2mac_dat_src_mask[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4141" *) sc2mac_dat_src_data75 : sc2mac_dat_data75_d1;
  assign _099_ = sc2mac_dat_src_mask[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4131" *) sc2mac_dat_src_data74 : sc2mac_dat_data74_d1;
  assign _098_ = sc2mac_dat_src_mask[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4121" *) sc2mac_dat_src_data73 : sc2mac_dat_data73_d1;
  assign _097_ = sc2mac_dat_src_mask[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4111" *) sc2mac_dat_src_data72 : sc2mac_dat_data72_d1;
  assign _096_ = sc2mac_dat_src_mask[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4101" *) sc2mac_dat_src_data71 : sc2mac_dat_data71_d1;
  assign _095_ = sc2mac_dat_src_mask[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4091" *) sc2mac_dat_src_data70 : sc2mac_dat_data70_d1;
  assign _093_ = sc2mac_dat_src_mask[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4081" *) sc2mac_dat_src_data69 : sc2mac_dat_data69_d1;
  assign _092_ = sc2mac_dat_src_mask[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4071" *) sc2mac_dat_src_data68 : sc2mac_dat_data68_d1;
  assign _091_ = sc2mac_dat_src_mask[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4061" *) sc2mac_dat_src_data67 : sc2mac_dat_data67_d1;
  assign _090_ = sc2mac_dat_src_mask[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4051" *) sc2mac_dat_src_data66 : sc2mac_dat_data66_d1;
  assign _089_ = sc2mac_dat_src_mask[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4041" *) sc2mac_dat_src_data65 : sc2mac_dat_data65_d1;
  assign _088_ = sc2mac_dat_src_mask[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4031" *) sc2mac_dat_src_data64 : sc2mac_dat_data64_d1;
  assign _087_ = sc2mac_dat_src_mask[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4021" *) sc2mac_dat_src_data63 : sc2mac_dat_data63_d1;
  assign _086_ = sc2mac_dat_src_mask[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4011" *) sc2mac_dat_src_data62 : sc2mac_dat_data62_d1;
  assign _085_ = sc2mac_dat_src_mask[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:4001" *) sc2mac_dat_src_data61 : sc2mac_dat_data61_d1;
  assign _084_ = sc2mac_dat_src_mask[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3991" *) sc2mac_dat_src_data60 : sc2mac_dat_data60_d1;
  assign _082_ = sc2mac_dat_src_mask[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3981" *) sc2mac_dat_src_data59 : sc2mac_dat_data59_d1;
  assign _081_ = sc2mac_dat_src_mask[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3971" *) sc2mac_dat_src_data58 : sc2mac_dat_data58_d1;
  assign _080_ = sc2mac_dat_src_mask[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3961" *) sc2mac_dat_src_data57 : sc2mac_dat_data57_d1;
  assign _079_ = sc2mac_dat_src_mask[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3951" *) sc2mac_dat_src_data56 : sc2mac_dat_data56_d1;
  assign _078_ = sc2mac_dat_src_mask[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3941" *) sc2mac_dat_src_data55 : sc2mac_dat_data55_d1;
  assign _077_ = sc2mac_dat_src_mask[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3931" *) sc2mac_dat_src_data54 : sc2mac_dat_data54_d1;
  assign _076_ = sc2mac_dat_src_mask[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3921" *) sc2mac_dat_src_data53 : sc2mac_dat_data53_d1;
  assign _075_ = sc2mac_dat_src_mask[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3911" *) sc2mac_dat_src_data52 : sc2mac_dat_data52_d1;
  assign _074_ = sc2mac_dat_src_mask[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3901" *) sc2mac_dat_src_data51 : sc2mac_dat_data51_d1;
  assign _073_ = sc2mac_dat_src_mask[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3891" *) sc2mac_dat_src_data50 : sc2mac_dat_data50_d1;
  assign _071_ = sc2mac_dat_src_mask[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3881" *) sc2mac_dat_src_data49 : sc2mac_dat_data49_d1;
  assign _070_ = sc2mac_dat_src_mask[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3871" *) sc2mac_dat_src_data48 : sc2mac_dat_data48_d1;
  assign _069_ = sc2mac_dat_src_mask[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3861" *) sc2mac_dat_src_data47 : sc2mac_dat_data47_d1;
  assign _068_ = sc2mac_dat_src_mask[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3851" *) sc2mac_dat_src_data46 : sc2mac_dat_data46_d1;
  assign _067_ = sc2mac_dat_src_mask[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3841" *) sc2mac_dat_src_data45 : sc2mac_dat_data45_d1;
  assign _066_ = sc2mac_dat_src_mask[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3831" *) sc2mac_dat_src_data44 : sc2mac_dat_data44_d1;
  assign _065_ = sc2mac_dat_src_mask[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3821" *) sc2mac_dat_src_data43 : sc2mac_dat_data43_d1;
  assign _064_ = sc2mac_dat_src_mask[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3811" *) sc2mac_dat_src_data42 : sc2mac_dat_data42_d1;
  assign _063_ = sc2mac_dat_src_mask[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3801" *) sc2mac_dat_src_data41 : sc2mac_dat_data41_d1;
  assign _062_ = sc2mac_dat_src_mask[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3791" *) sc2mac_dat_src_data40 : sc2mac_dat_data40_d1;
  assign _060_ = sc2mac_dat_src_mask[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3781" *) sc2mac_dat_src_data39 : sc2mac_dat_data39_d1;
  assign _059_ = sc2mac_dat_src_mask[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3771" *) sc2mac_dat_src_data38 : sc2mac_dat_data38_d1;
  assign _058_ = sc2mac_dat_src_mask[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3761" *) sc2mac_dat_src_data37 : sc2mac_dat_data37_d1;
  assign _057_ = sc2mac_dat_src_mask[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3751" *) sc2mac_dat_src_data36 : sc2mac_dat_data36_d1;
  assign _056_ = sc2mac_dat_src_mask[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3741" *) sc2mac_dat_src_data35 : sc2mac_dat_data35_d1;
  assign _055_ = sc2mac_dat_src_mask[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3731" *) sc2mac_dat_src_data34 : sc2mac_dat_data34_d1;
  assign _054_ = sc2mac_dat_src_mask[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3721" *) sc2mac_dat_src_data33 : sc2mac_dat_data33_d1;
  assign _053_ = sc2mac_dat_src_mask[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3711" *) sc2mac_dat_src_data32 : sc2mac_dat_data32_d1;
  assign _052_ = sc2mac_dat_src_mask[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3701" *) sc2mac_dat_src_data31 : sc2mac_dat_data31_d1;
  assign _051_ = sc2mac_dat_src_mask[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3691" *) sc2mac_dat_src_data30 : sc2mac_dat_data30_d1;
  assign _049_ = sc2mac_dat_src_mask[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3681" *) sc2mac_dat_src_data29 : sc2mac_dat_data29_d1;
  assign _048_ = sc2mac_dat_src_mask[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3671" *) sc2mac_dat_src_data28 : sc2mac_dat_data28_d1;
  assign _047_ = sc2mac_dat_src_mask[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3661" *) sc2mac_dat_src_data27 : sc2mac_dat_data27_d1;
  assign _046_ = sc2mac_dat_src_mask[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3651" *) sc2mac_dat_src_data26 : sc2mac_dat_data26_d1;
  assign _045_ = sc2mac_dat_src_mask[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3641" *) sc2mac_dat_src_data25 : sc2mac_dat_data25_d1;
  assign _044_ = sc2mac_dat_src_mask[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3631" *) sc2mac_dat_src_data24 : sc2mac_dat_data24_d1;
  assign _043_ = sc2mac_dat_src_mask[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3621" *) sc2mac_dat_src_data23 : sc2mac_dat_data23_d1;
  assign _042_ = sc2mac_dat_src_mask[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3611" *) sc2mac_dat_src_data22 : sc2mac_dat_data22_d1;
  assign _041_ = sc2mac_dat_src_mask[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3601" *) sc2mac_dat_src_data21 : sc2mac_dat_data21_d1;
  assign _040_ = sc2mac_dat_src_mask[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3591" *) sc2mac_dat_src_data20 : sc2mac_dat_data20_d1;
  assign _038_ = sc2mac_dat_src_mask[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3581" *) sc2mac_dat_src_data19 : sc2mac_dat_data19_d1;
  assign _037_ = sc2mac_dat_src_mask[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3571" *) sc2mac_dat_src_data18 : sc2mac_dat_data18_d1;
  assign _036_ = sc2mac_dat_src_mask[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3561" *) sc2mac_dat_src_data17 : sc2mac_dat_data17_d1;
  assign _035_ = sc2mac_dat_src_mask[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3551" *) sc2mac_dat_src_data16 : sc2mac_dat_data16_d1;
  assign _034_ = sc2mac_dat_src_mask[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3541" *) sc2mac_dat_src_data15 : sc2mac_dat_data15_d1;
  assign _033_ = sc2mac_dat_src_mask[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3531" *) sc2mac_dat_src_data14 : sc2mac_dat_data14_d1;
  assign _032_ = sc2mac_dat_src_mask[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3521" *) sc2mac_dat_src_data13 : sc2mac_dat_data13_d1;
  assign _031_ = sc2mac_dat_src_mask[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3511" *) sc2mac_dat_src_data12 : sc2mac_dat_data12_d1;
  assign _022_ = sc2mac_dat_src_mask[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3501" *) sc2mac_dat_src_data11 : sc2mac_dat_data11_d1;
  assign _011_ = sc2mac_dat_src_mask[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3491" *) sc2mac_dat_src_data10 : sc2mac_dat_data10_d1;
  assign _127_ = sc2mac_dat_src_mask[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3481" *) sc2mac_dat_src_data9 : sc2mac_dat_data9_d1;
  assign _116_ = sc2mac_dat_src_mask[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3471" *) sc2mac_dat_src_data8 : sc2mac_dat_data8_d1;
  assign _105_ = sc2mac_dat_src_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3461" *) sc2mac_dat_src_data7 : sc2mac_dat_data7_d1;
  assign _094_ = sc2mac_dat_src_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3451" *) sc2mac_dat_src_data6 : sc2mac_dat_data6_d1;
  assign _083_ = sc2mac_dat_src_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3441" *) sc2mac_dat_src_data5 : sc2mac_dat_data5_d1;
  assign _072_ = sc2mac_dat_src_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3431" *) sc2mac_dat_src_data4 : sc2mac_dat_data4_d1;
  assign _061_ = sc2mac_dat_src_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3421" *) sc2mac_dat_src_data3 : sc2mac_dat_data3_d1;
  assign _050_ = sc2mac_dat_src_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3411" *) sc2mac_dat_src_data2 : sc2mac_dat_data2_d1;
  assign _039_ = sc2mac_dat_src_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3401" *) sc2mac_dat_src_data1 : sc2mac_dat_data1_d1;
  assign _000_ = sc2mac_dat_src_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3391" *) sc2mac_dat_src_data0 : sc2mac_dat_data0_d1;
  assign _128_ = _261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3333" *) sc2mac_dat_src_mask : sc2mac_dat_mask_d1;
  assign _129_ = _261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3272" *) sc2mac_dat_src_pd : sc2mac_dat_pd_d1;
  assign _160_ = sc2mac_wt_src_mask[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3252" *) sc2mac_wt_src_data127 : sc2mac_wt_data127_d1;
  assign _159_ = sc2mac_wt_src_mask[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3242" *) sc2mac_wt_src_data126 : sc2mac_wt_data126_d1;
  assign _158_ = sc2mac_wt_src_mask[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3232" *) sc2mac_wt_src_data125 : sc2mac_wt_data125_d1;
  assign _157_ = sc2mac_wt_src_mask[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3222" *) sc2mac_wt_src_data124 : sc2mac_wt_data124_d1;
  assign _156_ = sc2mac_wt_src_mask[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3212" *) sc2mac_wt_src_data123 : sc2mac_wt_data123_d1;
  assign _155_ = sc2mac_wt_src_mask[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3202" *) sc2mac_wt_src_data122 : sc2mac_wt_data122_d1;
  assign _154_ = sc2mac_wt_src_mask[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3192" *) sc2mac_wt_src_data121 : sc2mac_wt_data121_d1;
  assign _153_ = sc2mac_wt_src_mask[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3182" *) sc2mac_wt_src_data120 : sc2mac_wt_data120_d1;
  assign _151_ = sc2mac_wt_src_mask[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3172" *) sc2mac_wt_src_data119 : sc2mac_wt_data119_d1;
  assign _150_ = sc2mac_wt_src_mask[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3162" *) sc2mac_wt_src_data118 : sc2mac_wt_data118_d1;
  assign _149_ = sc2mac_wt_src_mask[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3152" *) sc2mac_wt_src_data117 : sc2mac_wt_data117_d1;
  assign _148_ = sc2mac_wt_src_mask[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3142" *) sc2mac_wt_src_data116 : sc2mac_wt_data116_d1;
  assign _147_ = sc2mac_wt_src_mask[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3132" *) sc2mac_wt_src_data115 : sc2mac_wt_data115_d1;
  assign _146_ = sc2mac_wt_src_mask[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3122" *) sc2mac_wt_src_data114 : sc2mac_wt_data114_d1;
  assign _145_ = sc2mac_wt_src_mask[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3112" *) sc2mac_wt_src_data113 : sc2mac_wt_data113_d1;
  assign _144_ = sc2mac_wt_src_mask[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3102" *) sc2mac_wt_src_data112 : sc2mac_wt_data112_d1;
  assign _143_ = sc2mac_wt_src_mask[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3092" *) sc2mac_wt_src_data111 : sc2mac_wt_data111_d1;
  assign _142_ = sc2mac_wt_src_mask[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3082" *) sc2mac_wt_src_data110 : sc2mac_wt_data110_d1;
  assign _140_ = sc2mac_wt_src_mask[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3072" *) sc2mac_wt_src_data109 : sc2mac_wt_data109_d1;
  assign _139_ = sc2mac_wt_src_mask[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3062" *) sc2mac_wt_src_data108 : sc2mac_wt_data108_d1;
  assign _138_ = sc2mac_wt_src_mask[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3052" *) sc2mac_wt_src_data107 : sc2mac_wt_data107_d1;
  assign _137_ = sc2mac_wt_src_mask[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3042" *) sc2mac_wt_src_data106 : sc2mac_wt_data106_d1;
  assign _136_ = sc2mac_wt_src_mask[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3032" *) sc2mac_wt_src_data105 : sc2mac_wt_data105_d1;
  assign _135_ = sc2mac_wt_src_mask[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3022" *) sc2mac_wt_src_data104 : sc2mac_wt_data104_d1;
  assign _134_ = sc2mac_wt_src_mask[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3012" *) sc2mac_wt_src_data103 : sc2mac_wt_data103_d1;
  assign _133_ = sc2mac_wt_src_mask[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:3002" *) sc2mac_wt_src_data102 : sc2mac_wt_data102_d1;
  assign _132_ = sc2mac_wt_src_mask[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2992" *) sc2mac_wt_src_data101 : sc2mac_wt_data101_d1;
  assign _131_ = sc2mac_wt_src_mask[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2982" *) sc2mac_wt_src_data100 : sc2mac_wt_data100_d1;
  assign _256_ = sc2mac_wt_src_mask[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2972" *) sc2mac_wt_src_data99 : sc2mac_wt_data99_d1;
  assign _255_ = sc2mac_wt_src_mask[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2962" *) sc2mac_wt_src_data98 : sc2mac_wt_data98_d1;
  assign _254_ = sc2mac_wt_src_mask[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2952" *) sc2mac_wt_src_data97 : sc2mac_wt_data97_d1;
  assign _253_ = sc2mac_wt_src_mask[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2942" *) sc2mac_wt_src_data96 : sc2mac_wt_data96_d1;
  assign _252_ = sc2mac_wt_src_mask[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2932" *) sc2mac_wt_src_data95 : sc2mac_wt_data95_d1;
  assign _251_ = sc2mac_wt_src_mask[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2922" *) sc2mac_wt_src_data94 : sc2mac_wt_data94_d1;
  assign _250_ = sc2mac_wt_src_mask[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2912" *) sc2mac_wt_src_data93 : sc2mac_wt_data93_d1;
  assign _249_ = sc2mac_wt_src_mask[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2902" *) sc2mac_wt_src_data92 : sc2mac_wt_data92_d1;
  assign _248_ = sc2mac_wt_src_mask[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2892" *) sc2mac_wt_src_data91 : sc2mac_wt_data91_d1;
  assign _247_ = sc2mac_wt_src_mask[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2882" *) sc2mac_wt_src_data90 : sc2mac_wt_data90_d1;
  assign _245_ = sc2mac_wt_src_mask[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2872" *) sc2mac_wt_src_data89 : sc2mac_wt_data89_d1;
  assign _244_ = sc2mac_wt_src_mask[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2862" *) sc2mac_wt_src_data88 : sc2mac_wt_data88_d1;
  assign _243_ = sc2mac_wt_src_mask[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2852" *) sc2mac_wt_src_data87 : sc2mac_wt_data87_d1;
  assign _242_ = sc2mac_wt_src_mask[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2842" *) sc2mac_wt_src_data86 : sc2mac_wt_data86_d1;
  assign _241_ = sc2mac_wt_src_mask[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2832" *) sc2mac_wt_src_data85 : sc2mac_wt_data85_d1;
  assign _240_ = sc2mac_wt_src_mask[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2822" *) sc2mac_wt_src_data84 : sc2mac_wt_data84_d1;
  assign _239_ = sc2mac_wt_src_mask[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2812" *) sc2mac_wt_src_data83 : sc2mac_wt_data83_d1;
  assign _238_ = sc2mac_wt_src_mask[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2802" *) sc2mac_wt_src_data82 : sc2mac_wt_data82_d1;
  assign _237_ = sc2mac_wt_src_mask[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2792" *) sc2mac_wt_src_data81 : sc2mac_wt_data81_d1;
  assign _236_ = sc2mac_wt_src_mask[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2782" *) sc2mac_wt_src_data80 : sc2mac_wt_data80_d1;
  assign _234_ = sc2mac_wt_src_mask[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2772" *) sc2mac_wt_src_data79 : sc2mac_wt_data79_d1;
  assign _233_ = sc2mac_wt_src_mask[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2762" *) sc2mac_wt_src_data78 : sc2mac_wt_data78_d1;
  assign _232_ = sc2mac_wt_src_mask[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2752" *) sc2mac_wt_src_data77 : sc2mac_wt_data77_d1;
  assign _231_ = sc2mac_wt_src_mask[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2742" *) sc2mac_wt_src_data76 : sc2mac_wt_data76_d1;
  assign _230_ = sc2mac_wt_src_mask[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2732" *) sc2mac_wt_src_data75 : sc2mac_wt_data75_d1;
  assign _229_ = sc2mac_wt_src_mask[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2722" *) sc2mac_wt_src_data74 : sc2mac_wt_data74_d1;
  assign _228_ = sc2mac_wt_src_mask[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2712" *) sc2mac_wt_src_data73 : sc2mac_wt_data73_d1;
  assign _227_ = sc2mac_wt_src_mask[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2702" *) sc2mac_wt_src_data72 : sc2mac_wt_data72_d1;
  assign _226_ = sc2mac_wt_src_mask[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2692" *) sc2mac_wt_src_data71 : sc2mac_wt_data71_d1;
  assign _225_ = sc2mac_wt_src_mask[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2682" *) sc2mac_wt_src_data70 : sc2mac_wt_data70_d1;
  assign _223_ = sc2mac_wt_src_mask[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2672" *) sc2mac_wt_src_data69 : sc2mac_wt_data69_d1;
  assign _222_ = sc2mac_wt_src_mask[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2662" *) sc2mac_wt_src_data68 : sc2mac_wt_data68_d1;
  assign _221_ = sc2mac_wt_src_mask[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2652" *) sc2mac_wt_src_data67 : sc2mac_wt_data67_d1;
  assign _220_ = sc2mac_wt_src_mask[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2642" *) sc2mac_wt_src_data66 : sc2mac_wt_data66_d1;
  assign _219_ = sc2mac_wt_src_mask[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2632" *) sc2mac_wt_src_data65 : sc2mac_wt_data65_d1;
  assign _218_ = sc2mac_wt_src_mask[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2622" *) sc2mac_wt_src_data64 : sc2mac_wt_data64_d1;
  assign _217_ = sc2mac_wt_src_mask[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2612" *) sc2mac_wt_src_data63 : sc2mac_wt_data63_d1;
  assign _216_ = sc2mac_wt_src_mask[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2602" *) sc2mac_wt_src_data62 : sc2mac_wt_data62_d1;
  assign _215_ = sc2mac_wt_src_mask[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2592" *) sc2mac_wt_src_data61 : sc2mac_wt_data61_d1;
  assign _214_ = sc2mac_wt_src_mask[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2582" *) sc2mac_wt_src_data60 : sc2mac_wt_data60_d1;
  assign _212_ = sc2mac_wt_src_mask[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2572" *) sc2mac_wt_src_data59 : sc2mac_wt_data59_d1;
  assign _211_ = sc2mac_wt_src_mask[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2562" *) sc2mac_wt_src_data58 : sc2mac_wt_data58_d1;
  assign _210_ = sc2mac_wt_src_mask[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2552" *) sc2mac_wt_src_data57 : sc2mac_wt_data57_d1;
  assign _209_ = sc2mac_wt_src_mask[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2542" *) sc2mac_wt_src_data56 : sc2mac_wt_data56_d1;
  assign _208_ = sc2mac_wt_src_mask[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2532" *) sc2mac_wt_src_data55 : sc2mac_wt_data55_d1;
  assign _207_ = sc2mac_wt_src_mask[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2522" *) sc2mac_wt_src_data54 : sc2mac_wt_data54_d1;
  assign _206_ = sc2mac_wt_src_mask[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2512" *) sc2mac_wt_src_data53 : sc2mac_wt_data53_d1;
  assign _205_ = sc2mac_wt_src_mask[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2502" *) sc2mac_wt_src_data52 : sc2mac_wt_data52_d1;
  assign _204_ = sc2mac_wt_src_mask[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2492" *) sc2mac_wt_src_data51 : sc2mac_wt_data51_d1;
  assign _203_ = sc2mac_wt_src_mask[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2482" *) sc2mac_wt_src_data50 : sc2mac_wt_data50_d1;
  assign _201_ = sc2mac_wt_src_mask[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2472" *) sc2mac_wt_src_data49 : sc2mac_wt_data49_d1;
  assign _200_ = sc2mac_wt_src_mask[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2462" *) sc2mac_wt_src_data48 : sc2mac_wt_data48_d1;
  assign _199_ = sc2mac_wt_src_mask[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2452" *) sc2mac_wt_src_data47 : sc2mac_wt_data47_d1;
  assign _198_ = sc2mac_wt_src_mask[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2442" *) sc2mac_wt_src_data46 : sc2mac_wt_data46_d1;
  assign _197_ = sc2mac_wt_src_mask[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2432" *) sc2mac_wt_src_data45 : sc2mac_wt_data45_d1;
  assign _196_ = sc2mac_wt_src_mask[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2422" *) sc2mac_wt_src_data44 : sc2mac_wt_data44_d1;
  assign _195_ = sc2mac_wt_src_mask[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2412" *) sc2mac_wt_src_data43 : sc2mac_wt_data43_d1;
  assign _194_ = sc2mac_wt_src_mask[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2402" *) sc2mac_wt_src_data42 : sc2mac_wt_data42_d1;
  assign _193_ = sc2mac_wt_src_mask[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2392" *) sc2mac_wt_src_data41 : sc2mac_wt_data41_d1;
  assign _192_ = sc2mac_wt_src_mask[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2382" *) sc2mac_wt_src_data40 : sc2mac_wt_data40_d1;
  assign _190_ = sc2mac_wt_src_mask[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2372" *) sc2mac_wt_src_data39 : sc2mac_wt_data39_d1;
  assign _189_ = sc2mac_wt_src_mask[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2362" *) sc2mac_wt_src_data38 : sc2mac_wt_data38_d1;
  assign _188_ = sc2mac_wt_src_mask[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2352" *) sc2mac_wt_src_data37 : sc2mac_wt_data37_d1;
  assign _187_ = sc2mac_wt_src_mask[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2342" *) sc2mac_wt_src_data36 : sc2mac_wt_data36_d1;
  assign _186_ = sc2mac_wt_src_mask[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2332" *) sc2mac_wt_src_data35 : sc2mac_wt_data35_d1;
  assign _185_ = sc2mac_wt_src_mask[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2322" *) sc2mac_wt_src_data34 : sc2mac_wt_data34_d1;
  assign _184_ = sc2mac_wt_src_mask[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2312" *) sc2mac_wt_src_data33 : sc2mac_wt_data33_d1;
  assign _183_ = sc2mac_wt_src_mask[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2302" *) sc2mac_wt_src_data32 : sc2mac_wt_data32_d1;
  assign _182_ = sc2mac_wt_src_mask[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2292" *) sc2mac_wt_src_data31 : sc2mac_wt_data31_d1;
  assign _181_ = sc2mac_wt_src_mask[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2282" *) sc2mac_wt_src_data30 : sc2mac_wt_data30_d1;
  assign _179_ = sc2mac_wt_src_mask[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2272" *) sc2mac_wt_src_data29 : sc2mac_wt_data29_d1;
  assign _178_ = sc2mac_wt_src_mask[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2262" *) sc2mac_wt_src_data28 : sc2mac_wt_data28_d1;
  assign _177_ = sc2mac_wt_src_mask[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2252" *) sc2mac_wt_src_data27 : sc2mac_wt_data27_d1;
  assign _176_ = sc2mac_wt_src_mask[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2242" *) sc2mac_wt_src_data26 : sc2mac_wt_data26_d1;
  assign _175_ = sc2mac_wt_src_mask[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2232" *) sc2mac_wt_src_data25 : sc2mac_wt_data25_d1;
  assign _174_ = sc2mac_wt_src_mask[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2222" *) sc2mac_wt_src_data24 : sc2mac_wt_data24_d1;
  assign _173_ = sc2mac_wt_src_mask[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2212" *) sc2mac_wt_src_data23 : sc2mac_wt_data23_d1;
  assign _172_ = sc2mac_wt_src_mask[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2202" *) sc2mac_wt_src_data22 : sc2mac_wt_data22_d1;
  assign _171_ = sc2mac_wt_src_mask[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2192" *) sc2mac_wt_src_data21 : sc2mac_wt_data21_d1;
  assign _170_ = sc2mac_wt_src_mask[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2182" *) sc2mac_wt_src_data20 : sc2mac_wt_data20_d1;
  assign _168_ = sc2mac_wt_src_mask[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2172" *) sc2mac_wt_src_data19 : sc2mac_wt_data19_d1;
  assign _167_ = sc2mac_wt_src_mask[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2162" *) sc2mac_wt_src_data18 : sc2mac_wt_data18_d1;
  assign _166_ = sc2mac_wt_src_mask[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2152" *) sc2mac_wt_src_data17 : sc2mac_wt_data17_d1;
  assign _165_ = sc2mac_wt_src_mask[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2142" *) sc2mac_wt_src_data16 : sc2mac_wt_data16_d1;
  assign _164_ = sc2mac_wt_src_mask[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2132" *) sc2mac_wt_src_data15 : sc2mac_wt_data15_d1;
  assign _163_ = sc2mac_wt_src_mask[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2122" *) sc2mac_wt_src_data14 : sc2mac_wt_data14_d1;
  assign _162_ = sc2mac_wt_src_mask[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2112" *) sc2mac_wt_src_data13 : sc2mac_wt_data13_d1;
  assign _161_ = sc2mac_wt_src_mask[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2102" *) sc2mac_wt_src_data12 : sc2mac_wt_data12_d1;
  assign _152_ = sc2mac_wt_src_mask[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2092" *) sc2mac_wt_src_data11 : sc2mac_wt_data11_d1;
  assign _141_ = sc2mac_wt_src_mask[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2082" *) sc2mac_wt_src_data10 : sc2mac_wt_data10_d1;
  assign _257_ = sc2mac_wt_src_mask[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2072" *) sc2mac_wt_src_data9 : sc2mac_wt_data9_d1;
  assign _246_ = sc2mac_wt_src_mask[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2062" *) sc2mac_wt_src_data8 : sc2mac_wt_data8_d1;
  assign _235_ = sc2mac_wt_src_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2052" *) sc2mac_wt_src_data7 : sc2mac_wt_data7_d1;
  assign _224_ = sc2mac_wt_src_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2042" *) sc2mac_wt_src_data6 : sc2mac_wt_data6_d1;
  assign _213_ = sc2mac_wt_src_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2032" *) sc2mac_wt_src_data5 : sc2mac_wt_data5_d1;
  assign _202_ = sc2mac_wt_src_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2022" *) sc2mac_wt_src_data4 : sc2mac_wt_data4_d1;
  assign _191_ = sc2mac_wt_src_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2012" *) sc2mac_wt_src_data3 : sc2mac_wt_data3_d1;
  assign _180_ = sc2mac_wt_src_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:2002" *) sc2mac_wt_src_data2 : sc2mac_wt_data2_d1;
  assign _169_ = sc2mac_wt_src_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1992" *) sc2mac_wt_src_data1 : sc2mac_wt_data1_d1;
  assign _130_ = sc2mac_wt_src_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1982" *) sc2mac_wt_src_data0 : sc2mac_wt_data0_d1;
  assign _258_ = _260_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1924" *) sc2mac_wt_src_mask : sc2mac_wt_mask_d1;
  assign _259_ = _260_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/retiming/NV_NVDLA_RT_csc2cmac_b.v:1863" *) sc2mac_wt_src_sel : sc2mac_wt_sel_d1;
  assign sc2mac_dat_data0_d0 = sc2mac_dat_src_data0;
  assign sc2mac_dat_data100_d0 = sc2mac_dat_src_data100;
  assign sc2mac_dat_data101_d0 = sc2mac_dat_src_data101;
  assign sc2mac_dat_data102_d0 = sc2mac_dat_src_data102;
  assign sc2mac_dat_data103_d0 = sc2mac_dat_src_data103;
  assign sc2mac_dat_data104_d0 = sc2mac_dat_src_data104;
  assign sc2mac_dat_data105_d0 = sc2mac_dat_src_data105;
  assign sc2mac_dat_data106_d0 = sc2mac_dat_src_data106;
  assign sc2mac_dat_data107_d0 = sc2mac_dat_src_data107;
  assign sc2mac_dat_data108_d0 = sc2mac_dat_src_data108;
  assign sc2mac_dat_data109_d0 = sc2mac_dat_src_data109;
  assign sc2mac_dat_data10_d0 = sc2mac_dat_src_data10;
  assign sc2mac_dat_data110_d0 = sc2mac_dat_src_data110;
  assign sc2mac_dat_data111_d0 = sc2mac_dat_src_data111;
  assign sc2mac_dat_data112_d0 = sc2mac_dat_src_data112;
  assign sc2mac_dat_data113_d0 = sc2mac_dat_src_data113;
  assign sc2mac_dat_data114_d0 = sc2mac_dat_src_data114;
  assign sc2mac_dat_data115_d0 = sc2mac_dat_src_data115;
  assign sc2mac_dat_data116_d0 = sc2mac_dat_src_data116;
  assign sc2mac_dat_data117_d0 = sc2mac_dat_src_data117;
  assign sc2mac_dat_data118_d0 = sc2mac_dat_src_data118;
  assign sc2mac_dat_data119_d0 = sc2mac_dat_src_data119;
  assign sc2mac_dat_data11_d0 = sc2mac_dat_src_data11;
  assign sc2mac_dat_data120_d0 = sc2mac_dat_src_data120;
  assign sc2mac_dat_data121_d0 = sc2mac_dat_src_data121;
  assign sc2mac_dat_data122_d0 = sc2mac_dat_src_data122;
  assign sc2mac_dat_data123_d0 = sc2mac_dat_src_data123;
  assign sc2mac_dat_data124_d0 = sc2mac_dat_src_data124;
  assign sc2mac_dat_data125_d0 = sc2mac_dat_src_data125;
  assign sc2mac_dat_data126_d0 = sc2mac_dat_src_data126;
  assign sc2mac_dat_data127_d0 = sc2mac_dat_src_data127;
  assign sc2mac_dat_data12_d0 = sc2mac_dat_src_data12;
  assign sc2mac_dat_data13_d0 = sc2mac_dat_src_data13;
  assign sc2mac_dat_data14_d0 = sc2mac_dat_src_data14;
  assign sc2mac_dat_data15_d0 = sc2mac_dat_src_data15;
  assign sc2mac_dat_data16_d0 = sc2mac_dat_src_data16;
  assign sc2mac_dat_data17_d0 = sc2mac_dat_src_data17;
  assign sc2mac_dat_data18_d0 = sc2mac_dat_src_data18;
  assign sc2mac_dat_data19_d0 = sc2mac_dat_src_data19;
  assign sc2mac_dat_data1_d0 = sc2mac_dat_src_data1;
  assign sc2mac_dat_data20_d0 = sc2mac_dat_src_data20;
  assign sc2mac_dat_data21_d0 = sc2mac_dat_src_data21;
  assign sc2mac_dat_data22_d0 = sc2mac_dat_src_data22;
  assign sc2mac_dat_data23_d0 = sc2mac_dat_src_data23;
  assign sc2mac_dat_data24_d0 = sc2mac_dat_src_data24;
  assign sc2mac_dat_data25_d0 = sc2mac_dat_src_data25;
  assign sc2mac_dat_data26_d0 = sc2mac_dat_src_data26;
  assign sc2mac_dat_data27_d0 = sc2mac_dat_src_data27;
  assign sc2mac_dat_data28_d0 = sc2mac_dat_src_data28;
  assign sc2mac_dat_data29_d0 = sc2mac_dat_src_data29;
  assign sc2mac_dat_data2_d0 = sc2mac_dat_src_data2;
  assign sc2mac_dat_data30_d0 = sc2mac_dat_src_data30;
  assign sc2mac_dat_data31_d0 = sc2mac_dat_src_data31;
  assign sc2mac_dat_data32_d0 = sc2mac_dat_src_data32;
  assign sc2mac_dat_data33_d0 = sc2mac_dat_src_data33;
  assign sc2mac_dat_data34_d0 = sc2mac_dat_src_data34;
  assign sc2mac_dat_data35_d0 = sc2mac_dat_src_data35;
  assign sc2mac_dat_data36_d0 = sc2mac_dat_src_data36;
  assign sc2mac_dat_data37_d0 = sc2mac_dat_src_data37;
  assign sc2mac_dat_data38_d0 = sc2mac_dat_src_data38;
  assign sc2mac_dat_data39_d0 = sc2mac_dat_src_data39;
  assign sc2mac_dat_data3_d0 = sc2mac_dat_src_data3;
  assign sc2mac_dat_data40_d0 = sc2mac_dat_src_data40;
  assign sc2mac_dat_data41_d0 = sc2mac_dat_src_data41;
  assign sc2mac_dat_data42_d0 = sc2mac_dat_src_data42;
  assign sc2mac_dat_data43_d0 = sc2mac_dat_src_data43;
  assign sc2mac_dat_data44_d0 = sc2mac_dat_src_data44;
  assign sc2mac_dat_data45_d0 = sc2mac_dat_src_data45;
  assign sc2mac_dat_data46_d0 = sc2mac_dat_src_data46;
  assign sc2mac_dat_data47_d0 = sc2mac_dat_src_data47;
  assign sc2mac_dat_data48_d0 = sc2mac_dat_src_data48;
  assign sc2mac_dat_data49_d0 = sc2mac_dat_src_data49;
  assign sc2mac_dat_data4_d0 = sc2mac_dat_src_data4;
  assign sc2mac_dat_data50_d0 = sc2mac_dat_src_data50;
  assign sc2mac_dat_data51_d0 = sc2mac_dat_src_data51;
  assign sc2mac_dat_data52_d0 = sc2mac_dat_src_data52;
  assign sc2mac_dat_data53_d0 = sc2mac_dat_src_data53;
  assign sc2mac_dat_data54_d0 = sc2mac_dat_src_data54;
  assign sc2mac_dat_data55_d0 = sc2mac_dat_src_data55;
  assign sc2mac_dat_data56_d0 = sc2mac_dat_src_data56;
  assign sc2mac_dat_data57_d0 = sc2mac_dat_src_data57;
  assign sc2mac_dat_data58_d0 = sc2mac_dat_src_data58;
  assign sc2mac_dat_data59_d0 = sc2mac_dat_src_data59;
  assign sc2mac_dat_data5_d0 = sc2mac_dat_src_data5;
  assign sc2mac_dat_data60_d0 = sc2mac_dat_src_data60;
  assign sc2mac_dat_data61_d0 = sc2mac_dat_src_data61;
  assign sc2mac_dat_data62_d0 = sc2mac_dat_src_data62;
  assign sc2mac_dat_data63_d0 = sc2mac_dat_src_data63;
  assign sc2mac_dat_data64_d0 = sc2mac_dat_src_data64;
  assign sc2mac_dat_data65_d0 = sc2mac_dat_src_data65;
  assign sc2mac_dat_data66_d0 = sc2mac_dat_src_data66;
  assign sc2mac_dat_data67_d0 = sc2mac_dat_src_data67;
  assign sc2mac_dat_data68_d0 = sc2mac_dat_src_data68;
  assign sc2mac_dat_data69_d0 = sc2mac_dat_src_data69;
  assign sc2mac_dat_data6_d0 = sc2mac_dat_src_data6;
  assign sc2mac_dat_data70_d0 = sc2mac_dat_src_data70;
  assign sc2mac_dat_data71_d0 = sc2mac_dat_src_data71;
  assign sc2mac_dat_data72_d0 = sc2mac_dat_src_data72;
  assign sc2mac_dat_data73_d0 = sc2mac_dat_src_data73;
  assign sc2mac_dat_data74_d0 = sc2mac_dat_src_data74;
  assign sc2mac_dat_data75_d0 = sc2mac_dat_src_data75;
  assign sc2mac_dat_data76_d0 = sc2mac_dat_src_data76;
  assign sc2mac_dat_data77_d0 = sc2mac_dat_src_data77;
  assign sc2mac_dat_data78_d0 = sc2mac_dat_src_data78;
  assign sc2mac_dat_data79_d0 = sc2mac_dat_src_data79;
  assign sc2mac_dat_data7_d0 = sc2mac_dat_src_data7;
  assign sc2mac_dat_data80_d0 = sc2mac_dat_src_data80;
  assign sc2mac_dat_data81_d0 = sc2mac_dat_src_data81;
  assign sc2mac_dat_data82_d0 = sc2mac_dat_src_data82;
  assign sc2mac_dat_data83_d0 = sc2mac_dat_src_data83;
  assign sc2mac_dat_data84_d0 = sc2mac_dat_src_data84;
  assign sc2mac_dat_data85_d0 = sc2mac_dat_src_data85;
  assign sc2mac_dat_data86_d0 = sc2mac_dat_src_data86;
  assign sc2mac_dat_data87_d0 = sc2mac_dat_src_data87;
  assign sc2mac_dat_data88_d0 = sc2mac_dat_src_data88;
  assign sc2mac_dat_data89_d0 = sc2mac_dat_src_data89;
  assign sc2mac_dat_data8_d0 = sc2mac_dat_src_data8;
  assign sc2mac_dat_data90_d0 = sc2mac_dat_src_data90;
  assign sc2mac_dat_data91_d0 = sc2mac_dat_src_data91;
  assign sc2mac_dat_data92_d0 = sc2mac_dat_src_data92;
  assign sc2mac_dat_data93_d0 = sc2mac_dat_src_data93;
  assign sc2mac_dat_data94_d0 = sc2mac_dat_src_data94;
  assign sc2mac_dat_data95_d0 = sc2mac_dat_src_data95;
  assign sc2mac_dat_data96_d0 = sc2mac_dat_src_data96;
  assign sc2mac_dat_data97_d0 = sc2mac_dat_src_data97;
  assign sc2mac_dat_data98_d0 = sc2mac_dat_src_data98;
  assign sc2mac_dat_data99_d0 = sc2mac_dat_src_data99;
  assign sc2mac_dat_data9_d0 = sc2mac_dat_src_data9;
  assign sc2mac_dat_dst_data0 = sc2mac_dat_data0_d1;
  assign sc2mac_dat_dst_data1 = sc2mac_dat_data1_d1;
  assign sc2mac_dat_dst_data10 = sc2mac_dat_data10_d1;
  assign sc2mac_dat_dst_data100 = sc2mac_dat_data100_d1;
  assign sc2mac_dat_dst_data101 = sc2mac_dat_data101_d1;
  assign sc2mac_dat_dst_data102 = sc2mac_dat_data102_d1;
  assign sc2mac_dat_dst_data103 = sc2mac_dat_data103_d1;
  assign sc2mac_dat_dst_data104 = sc2mac_dat_data104_d1;
  assign sc2mac_dat_dst_data105 = sc2mac_dat_data105_d1;
  assign sc2mac_dat_dst_data106 = sc2mac_dat_data106_d1;
  assign sc2mac_dat_dst_data107 = sc2mac_dat_data107_d1;
  assign sc2mac_dat_dst_data108 = sc2mac_dat_data108_d1;
  assign sc2mac_dat_dst_data109 = sc2mac_dat_data109_d1;
  assign sc2mac_dat_dst_data11 = sc2mac_dat_data11_d1;
  assign sc2mac_dat_dst_data110 = sc2mac_dat_data110_d1;
  assign sc2mac_dat_dst_data111 = sc2mac_dat_data111_d1;
  assign sc2mac_dat_dst_data112 = sc2mac_dat_data112_d1;
  assign sc2mac_dat_dst_data113 = sc2mac_dat_data113_d1;
  assign sc2mac_dat_dst_data114 = sc2mac_dat_data114_d1;
  assign sc2mac_dat_dst_data115 = sc2mac_dat_data115_d1;
  assign sc2mac_dat_dst_data116 = sc2mac_dat_data116_d1;
  assign sc2mac_dat_dst_data117 = sc2mac_dat_data117_d1;
  assign sc2mac_dat_dst_data118 = sc2mac_dat_data118_d1;
  assign sc2mac_dat_dst_data119 = sc2mac_dat_data119_d1;
  assign sc2mac_dat_dst_data12 = sc2mac_dat_data12_d1;
  assign sc2mac_dat_dst_data120 = sc2mac_dat_data120_d1;
  assign sc2mac_dat_dst_data121 = sc2mac_dat_data121_d1;
  assign sc2mac_dat_dst_data122 = sc2mac_dat_data122_d1;
  assign sc2mac_dat_dst_data123 = sc2mac_dat_data123_d1;
  assign sc2mac_dat_dst_data124 = sc2mac_dat_data124_d1;
  assign sc2mac_dat_dst_data125 = sc2mac_dat_data125_d1;
  assign sc2mac_dat_dst_data126 = sc2mac_dat_data126_d1;
  assign sc2mac_dat_dst_data127 = sc2mac_dat_data127_d1;
  assign sc2mac_dat_dst_data13 = sc2mac_dat_data13_d1;
  assign sc2mac_dat_dst_data14 = sc2mac_dat_data14_d1;
  assign sc2mac_dat_dst_data15 = sc2mac_dat_data15_d1;
  assign sc2mac_dat_dst_data16 = sc2mac_dat_data16_d1;
  assign sc2mac_dat_dst_data17 = sc2mac_dat_data17_d1;
  assign sc2mac_dat_dst_data18 = sc2mac_dat_data18_d1;
  assign sc2mac_dat_dst_data19 = sc2mac_dat_data19_d1;
  assign sc2mac_dat_dst_data2 = sc2mac_dat_data2_d1;
  assign sc2mac_dat_dst_data20 = sc2mac_dat_data20_d1;
  assign sc2mac_dat_dst_data21 = sc2mac_dat_data21_d1;
  assign sc2mac_dat_dst_data22 = sc2mac_dat_data22_d1;
  assign sc2mac_dat_dst_data23 = sc2mac_dat_data23_d1;
  assign sc2mac_dat_dst_data24 = sc2mac_dat_data24_d1;
  assign sc2mac_dat_dst_data25 = sc2mac_dat_data25_d1;
  assign sc2mac_dat_dst_data26 = sc2mac_dat_data26_d1;
  assign sc2mac_dat_dst_data27 = sc2mac_dat_data27_d1;
  assign sc2mac_dat_dst_data28 = sc2mac_dat_data28_d1;
  assign sc2mac_dat_dst_data29 = sc2mac_dat_data29_d1;
  assign sc2mac_dat_dst_data3 = sc2mac_dat_data3_d1;
  assign sc2mac_dat_dst_data30 = sc2mac_dat_data30_d1;
  assign sc2mac_dat_dst_data31 = sc2mac_dat_data31_d1;
  assign sc2mac_dat_dst_data32 = sc2mac_dat_data32_d1;
  assign sc2mac_dat_dst_data33 = sc2mac_dat_data33_d1;
  assign sc2mac_dat_dst_data34 = sc2mac_dat_data34_d1;
  assign sc2mac_dat_dst_data35 = sc2mac_dat_data35_d1;
  assign sc2mac_dat_dst_data36 = sc2mac_dat_data36_d1;
  assign sc2mac_dat_dst_data37 = sc2mac_dat_data37_d1;
  assign sc2mac_dat_dst_data38 = sc2mac_dat_data38_d1;
  assign sc2mac_dat_dst_data39 = sc2mac_dat_data39_d1;
  assign sc2mac_dat_dst_data4 = sc2mac_dat_data4_d1;
  assign sc2mac_dat_dst_data40 = sc2mac_dat_data40_d1;
  assign sc2mac_dat_dst_data41 = sc2mac_dat_data41_d1;
  assign sc2mac_dat_dst_data42 = sc2mac_dat_data42_d1;
  assign sc2mac_dat_dst_data43 = sc2mac_dat_data43_d1;
  assign sc2mac_dat_dst_data44 = sc2mac_dat_data44_d1;
  assign sc2mac_dat_dst_data45 = sc2mac_dat_data45_d1;
  assign sc2mac_dat_dst_data46 = sc2mac_dat_data46_d1;
  assign sc2mac_dat_dst_data47 = sc2mac_dat_data47_d1;
  assign sc2mac_dat_dst_data48 = sc2mac_dat_data48_d1;
  assign sc2mac_dat_dst_data49 = sc2mac_dat_data49_d1;
  assign sc2mac_dat_dst_data5 = sc2mac_dat_data5_d1;
  assign sc2mac_dat_dst_data50 = sc2mac_dat_data50_d1;
  assign sc2mac_dat_dst_data51 = sc2mac_dat_data51_d1;
  assign sc2mac_dat_dst_data52 = sc2mac_dat_data52_d1;
  assign sc2mac_dat_dst_data53 = sc2mac_dat_data53_d1;
  assign sc2mac_dat_dst_data54 = sc2mac_dat_data54_d1;
  assign sc2mac_dat_dst_data55 = sc2mac_dat_data55_d1;
  assign sc2mac_dat_dst_data56 = sc2mac_dat_data56_d1;
  assign sc2mac_dat_dst_data57 = sc2mac_dat_data57_d1;
  assign sc2mac_dat_dst_data58 = sc2mac_dat_data58_d1;
  assign sc2mac_dat_dst_data59 = sc2mac_dat_data59_d1;
  assign sc2mac_dat_dst_data6 = sc2mac_dat_data6_d1;
  assign sc2mac_dat_dst_data60 = sc2mac_dat_data60_d1;
  assign sc2mac_dat_dst_data61 = sc2mac_dat_data61_d1;
  assign sc2mac_dat_dst_data62 = sc2mac_dat_data62_d1;
  assign sc2mac_dat_dst_data63 = sc2mac_dat_data63_d1;
  assign sc2mac_dat_dst_data64 = sc2mac_dat_data64_d1;
  assign sc2mac_dat_dst_data65 = sc2mac_dat_data65_d1;
  assign sc2mac_dat_dst_data66 = sc2mac_dat_data66_d1;
  assign sc2mac_dat_dst_data67 = sc2mac_dat_data67_d1;
  assign sc2mac_dat_dst_data68 = sc2mac_dat_data68_d1;
  assign sc2mac_dat_dst_data69 = sc2mac_dat_data69_d1;
  assign sc2mac_dat_dst_data7 = sc2mac_dat_data7_d1;
  assign sc2mac_dat_dst_data70 = sc2mac_dat_data70_d1;
  assign sc2mac_dat_dst_data71 = sc2mac_dat_data71_d1;
  assign sc2mac_dat_dst_data72 = sc2mac_dat_data72_d1;
  assign sc2mac_dat_dst_data73 = sc2mac_dat_data73_d1;
  assign sc2mac_dat_dst_data74 = sc2mac_dat_data74_d1;
  assign sc2mac_dat_dst_data75 = sc2mac_dat_data75_d1;
  assign sc2mac_dat_dst_data76 = sc2mac_dat_data76_d1;
  assign sc2mac_dat_dst_data77 = sc2mac_dat_data77_d1;
  assign sc2mac_dat_dst_data78 = sc2mac_dat_data78_d1;
  assign sc2mac_dat_dst_data79 = sc2mac_dat_data79_d1;
  assign sc2mac_dat_dst_data8 = sc2mac_dat_data8_d1;
  assign sc2mac_dat_dst_data80 = sc2mac_dat_data80_d1;
  assign sc2mac_dat_dst_data81 = sc2mac_dat_data81_d1;
  assign sc2mac_dat_dst_data82 = sc2mac_dat_data82_d1;
  assign sc2mac_dat_dst_data83 = sc2mac_dat_data83_d1;
  assign sc2mac_dat_dst_data84 = sc2mac_dat_data84_d1;
  assign sc2mac_dat_dst_data85 = sc2mac_dat_data85_d1;
  assign sc2mac_dat_dst_data86 = sc2mac_dat_data86_d1;
  assign sc2mac_dat_dst_data87 = sc2mac_dat_data87_d1;
  assign sc2mac_dat_dst_data88 = sc2mac_dat_data88_d1;
  assign sc2mac_dat_dst_data89 = sc2mac_dat_data89_d1;
  assign sc2mac_dat_dst_data9 = sc2mac_dat_data9_d1;
  assign sc2mac_dat_dst_data90 = sc2mac_dat_data90_d1;
  assign sc2mac_dat_dst_data91 = sc2mac_dat_data91_d1;
  assign sc2mac_dat_dst_data92 = sc2mac_dat_data92_d1;
  assign sc2mac_dat_dst_data93 = sc2mac_dat_data93_d1;
  assign sc2mac_dat_dst_data94 = sc2mac_dat_data94_d1;
  assign sc2mac_dat_dst_data95 = sc2mac_dat_data95_d1;
  assign sc2mac_dat_dst_data96 = sc2mac_dat_data96_d1;
  assign sc2mac_dat_dst_data97 = sc2mac_dat_data97_d1;
  assign sc2mac_dat_dst_data98 = sc2mac_dat_data98_d1;
  assign sc2mac_dat_dst_data99 = sc2mac_dat_data99_d1;
  assign sc2mac_dat_dst_mask = sc2mac_dat_mask_d1;
  assign sc2mac_dat_dst_pd = sc2mac_dat_pd_d1;
  assign sc2mac_dat_dst_pvld = sc2mac_dat_pvld_d1;
  assign sc2mac_dat_mask_d0 = sc2mac_dat_src_mask;
  assign sc2mac_dat_pd_d0 = sc2mac_dat_src_pd;
  assign sc2mac_dat_pvld_d0 = sc2mac_dat_src_pvld;
  assign sc2mac_wt_data0_d0 = sc2mac_wt_src_data0;
  assign sc2mac_wt_data100_d0 = sc2mac_wt_src_data100;
  assign sc2mac_wt_data101_d0 = sc2mac_wt_src_data101;
  assign sc2mac_wt_data102_d0 = sc2mac_wt_src_data102;
  assign sc2mac_wt_data103_d0 = sc2mac_wt_src_data103;
  assign sc2mac_wt_data104_d0 = sc2mac_wt_src_data104;
  assign sc2mac_wt_data105_d0 = sc2mac_wt_src_data105;
  assign sc2mac_wt_data106_d0 = sc2mac_wt_src_data106;
  assign sc2mac_wt_data107_d0 = sc2mac_wt_src_data107;
  assign sc2mac_wt_data108_d0 = sc2mac_wt_src_data108;
  assign sc2mac_wt_data109_d0 = sc2mac_wt_src_data109;
  assign sc2mac_wt_data10_d0 = sc2mac_wt_src_data10;
  assign sc2mac_wt_data110_d0 = sc2mac_wt_src_data110;
  assign sc2mac_wt_data111_d0 = sc2mac_wt_src_data111;
  assign sc2mac_wt_data112_d0 = sc2mac_wt_src_data112;
  assign sc2mac_wt_data113_d0 = sc2mac_wt_src_data113;
  assign sc2mac_wt_data114_d0 = sc2mac_wt_src_data114;
  assign sc2mac_wt_data115_d0 = sc2mac_wt_src_data115;
  assign sc2mac_wt_data116_d0 = sc2mac_wt_src_data116;
  assign sc2mac_wt_data117_d0 = sc2mac_wt_src_data117;
  assign sc2mac_wt_data118_d0 = sc2mac_wt_src_data118;
  assign sc2mac_wt_data119_d0 = sc2mac_wt_src_data119;
  assign sc2mac_wt_data11_d0 = sc2mac_wt_src_data11;
  assign sc2mac_wt_data120_d0 = sc2mac_wt_src_data120;
  assign sc2mac_wt_data121_d0 = sc2mac_wt_src_data121;
  assign sc2mac_wt_data122_d0 = sc2mac_wt_src_data122;
  assign sc2mac_wt_data123_d0 = sc2mac_wt_src_data123;
  assign sc2mac_wt_data124_d0 = sc2mac_wt_src_data124;
  assign sc2mac_wt_data125_d0 = sc2mac_wt_src_data125;
  assign sc2mac_wt_data126_d0 = sc2mac_wt_src_data126;
  assign sc2mac_wt_data127_d0 = sc2mac_wt_src_data127;
  assign sc2mac_wt_data12_d0 = sc2mac_wt_src_data12;
  assign sc2mac_wt_data13_d0 = sc2mac_wt_src_data13;
  assign sc2mac_wt_data14_d0 = sc2mac_wt_src_data14;
  assign sc2mac_wt_data15_d0 = sc2mac_wt_src_data15;
  assign sc2mac_wt_data16_d0 = sc2mac_wt_src_data16;
  assign sc2mac_wt_data17_d0 = sc2mac_wt_src_data17;
  assign sc2mac_wt_data18_d0 = sc2mac_wt_src_data18;
  assign sc2mac_wt_data19_d0 = sc2mac_wt_src_data19;
  assign sc2mac_wt_data1_d0 = sc2mac_wt_src_data1;
  assign sc2mac_wt_data20_d0 = sc2mac_wt_src_data20;
  assign sc2mac_wt_data21_d0 = sc2mac_wt_src_data21;
  assign sc2mac_wt_data22_d0 = sc2mac_wt_src_data22;
  assign sc2mac_wt_data23_d0 = sc2mac_wt_src_data23;
  assign sc2mac_wt_data24_d0 = sc2mac_wt_src_data24;
  assign sc2mac_wt_data25_d0 = sc2mac_wt_src_data25;
  assign sc2mac_wt_data26_d0 = sc2mac_wt_src_data26;
  assign sc2mac_wt_data27_d0 = sc2mac_wt_src_data27;
  assign sc2mac_wt_data28_d0 = sc2mac_wt_src_data28;
  assign sc2mac_wt_data29_d0 = sc2mac_wt_src_data29;
  assign sc2mac_wt_data2_d0 = sc2mac_wt_src_data2;
  assign sc2mac_wt_data30_d0 = sc2mac_wt_src_data30;
  assign sc2mac_wt_data31_d0 = sc2mac_wt_src_data31;
  assign sc2mac_wt_data32_d0 = sc2mac_wt_src_data32;
  assign sc2mac_wt_data33_d0 = sc2mac_wt_src_data33;
  assign sc2mac_wt_data34_d0 = sc2mac_wt_src_data34;
  assign sc2mac_wt_data35_d0 = sc2mac_wt_src_data35;
  assign sc2mac_wt_data36_d0 = sc2mac_wt_src_data36;
  assign sc2mac_wt_data37_d0 = sc2mac_wt_src_data37;
  assign sc2mac_wt_data38_d0 = sc2mac_wt_src_data38;
  assign sc2mac_wt_data39_d0 = sc2mac_wt_src_data39;
  assign sc2mac_wt_data3_d0 = sc2mac_wt_src_data3;
  assign sc2mac_wt_data40_d0 = sc2mac_wt_src_data40;
  assign sc2mac_wt_data41_d0 = sc2mac_wt_src_data41;
  assign sc2mac_wt_data42_d0 = sc2mac_wt_src_data42;
  assign sc2mac_wt_data43_d0 = sc2mac_wt_src_data43;
  assign sc2mac_wt_data44_d0 = sc2mac_wt_src_data44;
  assign sc2mac_wt_data45_d0 = sc2mac_wt_src_data45;
  assign sc2mac_wt_data46_d0 = sc2mac_wt_src_data46;
  assign sc2mac_wt_data47_d0 = sc2mac_wt_src_data47;
  assign sc2mac_wt_data48_d0 = sc2mac_wt_src_data48;
  assign sc2mac_wt_data49_d0 = sc2mac_wt_src_data49;
  assign sc2mac_wt_data4_d0 = sc2mac_wt_src_data4;
  assign sc2mac_wt_data50_d0 = sc2mac_wt_src_data50;
  assign sc2mac_wt_data51_d0 = sc2mac_wt_src_data51;
  assign sc2mac_wt_data52_d0 = sc2mac_wt_src_data52;
  assign sc2mac_wt_data53_d0 = sc2mac_wt_src_data53;
  assign sc2mac_wt_data54_d0 = sc2mac_wt_src_data54;
  assign sc2mac_wt_data55_d0 = sc2mac_wt_src_data55;
  assign sc2mac_wt_data56_d0 = sc2mac_wt_src_data56;
  assign sc2mac_wt_data57_d0 = sc2mac_wt_src_data57;
  assign sc2mac_wt_data58_d0 = sc2mac_wt_src_data58;
  assign sc2mac_wt_data59_d0 = sc2mac_wt_src_data59;
  assign sc2mac_wt_data5_d0 = sc2mac_wt_src_data5;
  assign sc2mac_wt_data60_d0 = sc2mac_wt_src_data60;
  assign sc2mac_wt_data61_d0 = sc2mac_wt_src_data61;
  assign sc2mac_wt_data62_d0 = sc2mac_wt_src_data62;
  assign sc2mac_wt_data63_d0 = sc2mac_wt_src_data63;
  assign sc2mac_wt_data64_d0 = sc2mac_wt_src_data64;
  assign sc2mac_wt_data65_d0 = sc2mac_wt_src_data65;
  assign sc2mac_wt_data66_d0 = sc2mac_wt_src_data66;
  assign sc2mac_wt_data67_d0 = sc2mac_wt_src_data67;
  assign sc2mac_wt_data68_d0 = sc2mac_wt_src_data68;
  assign sc2mac_wt_data69_d0 = sc2mac_wt_src_data69;
  assign sc2mac_wt_data6_d0 = sc2mac_wt_src_data6;
  assign sc2mac_wt_data70_d0 = sc2mac_wt_src_data70;
  assign sc2mac_wt_data71_d0 = sc2mac_wt_src_data71;
  assign sc2mac_wt_data72_d0 = sc2mac_wt_src_data72;
  assign sc2mac_wt_data73_d0 = sc2mac_wt_src_data73;
  assign sc2mac_wt_data74_d0 = sc2mac_wt_src_data74;
  assign sc2mac_wt_data75_d0 = sc2mac_wt_src_data75;
  assign sc2mac_wt_data76_d0 = sc2mac_wt_src_data76;
  assign sc2mac_wt_data77_d0 = sc2mac_wt_src_data77;
  assign sc2mac_wt_data78_d0 = sc2mac_wt_src_data78;
  assign sc2mac_wt_data79_d0 = sc2mac_wt_src_data79;
  assign sc2mac_wt_data7_d0 = sc2mac_wt_src_data7;
  assign sc2mac_wt_data80_d0 = sc2mac_wt_src_data80;
  assign sc2mac_wt_data81_d0 = sc2mac_wt_src_data81;
  assign sc2mac_wt_data82_d0 = sc2mac_wt_src_data82;
  assign sc2mac_wt_data83_d0 = sc2mac_wt_src_data83;
  assign sc2mac_wt_data84_d0 = sc2mac_wt_src_data84;
  assign sc2mac_wt_data85_d0 = sc2mac_wt_src_data85;
  assign sc2mac_wt_data86_d0 = sc2mac_wt_src_data86;
  assign sc2mac_wt_data87_d0 = sc2mac_wt_src_data87;
  assign sc2mac_wt_data88_d0 = sc2mac_wt_src_data88;
  assign sc2mac_wt_data89_d0 = sc2mac_wt_src_data89;
  assign sc2mac_wt_data8_d0 = sc2mac_wt_src_data8;
  assign sc2mac_wt_data90_d0 = sc2mac_wt_src_data90;
  assign sc2mac_wt_data91_d0 = sc2mac_wt_src_data91;
  assign sc2mac_wt_data92_d0 = sc2mac_wt_src_data92;
  assign sc2mac_wt_data93_d0 = sc2mac_wt_src_data93;
  assign sc2mac_wt_data94_d0 = sc2mac_wt_src_data94;
  assign sc2mac_wt_data95_d0 = sc2mac_wt_src_data95;
  assign sc2mac_wt_data96_d0 = sc2mac_wt_src_data96;
  assign sc2mac_wt_data97_d0 = sc2mac_wt_src_data97;
  assign sc2mac_wt_data98_d0 = sc2mac_wt_src_data98;
  assign sc2mac_wt_data99_d0 = sc2mac_wt_src_data99;
  assign sc2mac_wt_data9_d0 = sc2mac_wt_src_data9;
  assign sc2mac_wt_dst_data0 = sc2mac_wt_data0_d1;
  assign sc2mac_wt_dst_data1 = sc2mac_wt_data1_d1;
  assign sc2mac_wt_dst_data10 = sc2mac_wt_data10_d1;
  assign sc2mac_wt_dst_data100 = sc2mac_wt_data100_d1;
  assign sc2mac_wt_dst_data101 = sc2mac_wt_data101_d1;
  assign sc2mac_wt_dst_data102 = sc2mac_wt_data102_d1;
  assign sc2mac_wt_dst_data103 = sc2mac_wt_data103_d1;
  assign sc2mac_wt_dst_data104 = sc2mac_wt_data104_d1;
  assign sc2mac_wt_dst_data105 = sc2mac_wt_data105_d1;
  assign sc2mac_wt_dst_data106 = sc2mac_wt_data106_d1;
  assign sc2mac_wt_dst_data107 = sc2mac_wt_data107_d1;
  assign sc2mac_wt_dst_data108 = sc2mac_wt_data108_d1;
  assign sc2mac_wt_dst_data109 = sc2mac_wt_data109_d1;
  assign sc2mac_wt_dst_data11 = sc2mac_wt_data11_d1;
  assign sc2mac_wt_dst_data110 = sc2mac_wt_data110_d1;
  assign sc2mac_wt_dst_data111 = sc2mac_wt_data111_d1;
  assign sc2mac_wt_dst_data112 = sc2mac_wt_data112_d1;
  assign sc2mac_wt_dst_data113 = sc2mac_wt_data113_d1;
  assign sc2mac_wt_dst_data114 = sc2mac_wt_data114_d1;
  assign sc2mac_wt_dst_data115 = sc2mac_wt_data115_d1;
  assign sc2mac_wt_dst_data116 = sc2mac_wt_data116_d1;
  assign sc2mac_wt_dst_data117 = sc2mac_wt_data117_d1;
  assign sc2mac_wt_dst_data118 = sc2mac_wt_data118_d1;
  assign sc2mac_wt_dst_data119 = sc2mac_wt_data119_d1;
  assign sc2mac_wt_dst_data12 = sc2mac_wt_data12_d1;
  assign sc2mac_wt_dst_data120 = sc2mac_wt_data120_d1;
  assign sc2mac_wt_dst_data121 = sc2mac_wt_data121_d1;
  assign sc2mac_wt_dst_data122 = sc2mac_wt_data122_d1;
  assign sc2mac_wt_dst_data123 = sc2mac_wt_data123_d1;
  assign sc2mac_wt_dst_data124 = sc2mac_wt_data124_d1;
  assign sc2mac_wt_dst_data125 = sc2mac_wt_data125_d1;
  assign sc2mac_wt_dst_data126 = sc2mac_wt_data126_d1;
  assign sc2mac_wt_dst_data127 = sc2mac_wt_data127_d1;
  assign sc2mac_wt_dst_data13 = sc2mac_wt_data13_d1;
  assign sc2mac_wt_dst_data14 = sc2mac_wt_data14_d1;
  assign sc2mac_wt_dst_data15 = sc2mac_wt_data15_d1;
  assign sc2mac_wt_dst_data16 = sc2mac_wt_data16_d1;
  assign sc2mac_wt_dst_data17 = sc2mac_wt_data17_d1;
  assign sc2mac_wt_dst_data18 = sc2mac_wt_data18_d1;
  assign sc2mac_wt_dst_data19 = sc2mac_wt_data19_d1;
  assign sc2mac_wt_dst_data2 = sc2mac_wt_data2_d1;
  assign sc2mac_wt_dst_data20 = sc2mac_wt_data20_d1;
  assign sc2mac_wt_dst_data21 = sc2mac_wt_data21_d1;
  assign sc2mac_wt_dst_data22 = sc2mac_wt_data22_d1;
  assign sc2mac_wt_dst_data23 = sc2mac_wt_data23_d1;
  assign sc2mac_wt_dst_data24 = sc2mac_wt_data24_d1;
  assign sc2mac_wt_dst_data25 = sc2mac_wt_data25_d1;
  assign sc2mac_wt_dst_data26 = sc2mac_wt_data26_d1;
  assign sc2mac_wt_dst_data27 = sc2mac_wt_data27_d1;
  assign sc2mac_wt_dst_data28 = sc2mac_wt_data28_d1;
  assign sc2mac_wt_dst_data29 = sc2mac_wt_data29_d1;
  assign sc2mac_wt_dst_data3 = sc2mac_wt_data3_d1;
  assign sc2mac_wt_dst_data30 = sc2mac_wt_data30_d1;
  assign sc2mac_wt_dst_data31 = sc2mac_wt_data31_d1;
  assign sc2mac_wt_dst_data32 = sc2mac_wt_data32_d1;
  assign sc2mac_wt_dst_data33 = sc2mac_wt_data33_d1;
  assign sc2mac_wt_dst_data34 = sc2mac_wt_data34_d1;
  assign sc2mac_wt_dst_data35 = sc2mac_wt_data35_d1;
  assign sc2mac_wt_dst_data36 = sc2mac_wt_data36_d1;
  assign sc2mac_wt_dst_data37 = sc2mac_wt_data37_d1;
  assign sc2mac_wt_dst_data38 = sc2mac_wt_data38_d1;
  assign sc2mac_wt_dst_data39 = sc2mac_wt_data39_d1;
  assign sc2mac_wt_dst_data4 = sc2mac_wt_data4_d1;
  assign sc2mac_wt_dst_data40 = sc2mac_wt_data40_d1;
  assign sc2mac_wt_dst_data41 = sc2mac_wt_data41_d1;
  assign sc2mac_wt_dst_data42 = sc2mac_wt_data42_d1;
  assign sc2mac_wt_dst_data43 = sc2mac_wt_data43_d1;
  assign sc2mac_wt_dst_data44 = sc2mac_wt_data44_d1;
  assign sc2mac_wt_dst_data45 = sc2mac_wt_data45_d1;
  assign sc2mac_wt_dst_data46 = sc2mac_wt_data46_d1;
  assign sc2mac_wt_dst_data47 = sc2mac_wt_data47_d1;
  assign sc2mac_wt_dst_data48 = sc2mac_wt_data48_d1;
  assign sc2mac_wt_dst_data49 = sc2mac_wt_data49_d1;
  assign sc2mac_wt_dst_data5 = sc2mac_wt_data5_d1;
  assign sc2mac_wt_dst_data50 = sc2mac_wt_data50_d1;
  assign sc2mac_wt_dst_data51 = sc2mac_wt_data51_d1;
  assign sc2mac_wt_dst_data52 = sc2mac_wt_data52_d1;
  assign sc2mac_wt_dst_data53 = sc2mac_wt_data53_d1;
  assign sc2mac_wt_dst_data54 = sc2mac_wt_data54_d1;
  assign sc2mac_wt_dst_data55 = sc2mac_wt_data55_d1;
  assign sc2mac_wt_dst_data56 = sc2mac_wt_data56_d1;
  assign sc2mac_wt_dst_data57 = sc2mac_wt_data57_d1;
  assign sc2mac_wt_dst_data58 = sc2mac_wt_data58_d1;
  assign sc2mac_wt_dst_data59 = sc2mac_wt_data59_d1;
  assign sc2mac_wt_dst_data6 = sc2mac_wt_data6_d1;
  assign sc2mac_wt_dst_data60 = sc2mac_wt_data60_d1;
  assign sc2mac_wt_dst_data61 = sc2mac_wt_data61_d1;
  assign sc2mac_wt_dst_data62 = sc2mac_wt_data62_d1;
  assign sc2mac_wt_dst_data63 = sc2mac_wt_data63_d1;
  assign sc2mac_wt_dst_data64 = sc2mac_wt_data64_d1;
  assign sc2mac_wt_dst_data65 = sc2mac_wt_data65_d1;
  assign sc2mac_wt_dst_data66 = sc2mac_wt_data66_d1;
  assign sc2mac_wt_dst_data67 = sc2mac_wt_data67_d1;
  assign sc2mac_wt_dst_data68 = sc2mac_wt_data68_d1;
  assign sc2mac_wt_dst_data69 = sc2mac_wt_data69_d1;
  assign sc2mac_wt_dst_data7 = sc2mac_wt_data7_d1;
  assign sc2mac_wt_dst_data70 = sc2mac_wt_data70_d1;
  assign sc2mac_wt_dst_data71 = sc2mac_wt_data71_d1;
  assign sc2mac_wt_dst_data72 = sc2mac_wt_data72_d1;
  assign sc2mac_wt_dst_data73 = sc2mac_wt_data73_d1;
  assign sc2mac_wt_dst_data74 = sc2mac_wt_data74_d1;
  assign sc2mac_wt_dst_data75 = sc2mac_wt_data75_d1;
  assign sc2mac_wt_dst_data76 = sc2mac_wt_data76_d1;
  assign sc2mac_wt_dst_data77 = sc2mac_wt_data77_d1;
  assign sc2mac_wt_dst_data78 = sc2mac_wt_data78_d1;
  assign sc2mac_wt_dst_data79 = sc2mac_wt_data79_d1;
  assign sc2mac_wt_dst_data8 = sc2mac_wt_data8_d1;
  assign sc2mac_wt_dst_data80 = sc2mac_wt_data80_d1;
  assign sc2mac_wt_dst_data81 = sc2mac_wt_data81_d1;
  assign sc2mac_wt_dst_data82 = sc2mac_wt_data82_d1;
  assign sc2mac_wt_dst_data83 = sc2mac_wt_data83_d1;
  assign sc2mac_wt_dst_data84 = sc2mac_wt_data84_d1;
  assign sc2mac_wt_dst_data85 = sc2mac_wt_data85_d1;
  assign sc2mac_wt_dst_data86 = sc2mac_wt_data86_d1;
  assign sc2mac_wt_dst_data87 = sc2mac_wt_data87_d1;
  assign sc2mac_wt_dst_data88 = sc2mac_wt_data88_d1;
  assign sc2mac_wt_dst_data89 = sc2mac_wt_data89_d1;
  assign sc2mac_wt_dst_data9 = sc2mac_wt_data9_d1;
  assign sc2mac_wt_dst_data90 = sc2mac_wt_data90_d1;
  assign sc2mac_wt_dst_data91 = sc2mac_wt_data91_d1;
  assign sc2mac_wt_dst_data92 = sc2mac_wt_data92_d1;
  assign sc2mac_wt_dst_data93 = sc2mac_wt_data93_d1;
  assign sc2mac_wt_dst_data94 = sc2mac_wt_data94_d1;
  assign sc2mac_wt_dst_data95 = sc2mac_wt_data95_d1;
  assign sc2mac_wt_dst_data96 = sc2mac_wt_data96_d1;
  assign sc2mac_wt_dst_data97 = sc2mac_wt_data97_d1;
  assign sc2mac_wt_dst_data98 = sc2mac_wt_data98_d1;
  assign sc2mac_wt_dst_data99 = sc2mac_wt_data99_d1;
  assign sc2mac_wt_dst_mask = sc2mac_wt_mask_d1;
  assign sc2mac_wt_dst_pvld = sc2mac_wt_pvld_d1;
  assign sc2mac_wt_dst_sel = sc2mac_wt_sel_d1;
  assign sc2mac_wt_mask_d0 = sc2mac_wt_src_mask;
  assign sc2mac_wt_pvld_d0 = sc2mac_wt_src_pvld;
  assign sc2mac_wt_sel_d0 = sc2mac_wt_src_sel;
endmodule
