module NV_NVDLA_PDP_CORE_cal2d(nvdla_core_clk, nvdla_core_rstn, nvdla_op_gated_clk_fp16, padding_v_cfg, pdp_dp2wdma_ready, pdp_op_start, pooling1d_pd, pooling1d_pvld, pooling_channel_cfg, pooling_out_fwidth_cfg, pooling_out_lwidth_cfg, pooling_out_mwidth_cfg, pooling_size_v_cfg, pooling_splitw_num_cfg, pooling_stride_v_cfg, pooling_type_cfg, pwrbus_ram_pd, reg2dp_cube_in_height, reg2dp_cube_out_width, reg2dp_fp16_en, reg2dp_input_data, reg2dp_int16_en, reg2dp_int8_en, reg2dp_kernel_height, reg2dp_kernel_width, reg2dp_pad_bottom_cfg, reg2dp_pad_top, reg2dp_pad_value_1x_cfg, reg2dp_pad_value_2x_cfg, reg2dp_pad_value_3x_cfg, reg2dp_pad_value_4x_cfg, reg2dp_pad_value_5x_cfg, reg2dp_pad_value_6x_cfg, reg2dp_pad_value_7x_cfg, reg2dp_partial_width_out_first, reg2dp_partial_width_out_last, reg2dp_partial_width_out_mid, reg2dp_recip_height_cfg, reg2dp_recip_width_cfg, pdp_dp2wdma_pd, pdp_dp2wdma_valid, pooling1d_prdy);
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0000_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0001_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0002_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0003_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0004_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0005_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0006_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0007_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0008_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0009_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0010_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0011_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0012_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0013_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0014_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0015_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0016_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0017_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0018_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0019_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0020_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0021_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0022_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0023_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0024_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0025_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0026_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0027_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0028_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0029_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0030_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0031_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0032_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0033_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0034_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0035_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0036_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0037_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0038_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0039_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0040_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0041_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0042_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0043_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0044_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0045_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0046_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0047_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0048_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0049_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0050_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0051_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0052_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0053_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0054_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0055_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0056_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0057_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0058_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0059_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0060_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0061_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0062_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0063_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0064_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0065_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0066_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0067_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0068_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0069_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0070_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0071_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0072_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0073_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0074_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0075_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0076_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0077_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0078_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0079_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0080_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0081_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0082_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0083_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0084_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0085_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0086_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0087_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0088_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0089_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0090_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0091_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0092_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0093_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0094_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0095_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0096_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0097_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0098_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0099_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0100_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0101_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0102_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0103_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0104_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0105_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0106_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0107_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0108_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0109_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0110_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0111_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0112_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0113_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0114_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0115_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0116_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0117_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0118_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0119_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0120_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0121_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0122_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0123_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0124_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0125_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0126_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0127_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0128_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0129_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0130_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0131_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0132_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0133_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0134_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0135_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0136_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0137_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0138_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0139_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0140_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0141_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0142_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0143_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0144_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0145_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0146_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0147_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0148_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0149_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0150_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0151_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0152_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0153_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0154_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0155_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0156_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0157_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0158_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0159_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0160_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0161_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0162_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0163_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0164_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0165_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0166_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0167_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0168_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0169_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0170_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0171_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0172_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0173_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0174_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0175_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0176_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0177_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0178_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0179_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0180_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0181_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0182_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0183_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0184_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0185_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0186_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0187_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0188_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0189_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0190_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0191_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0192_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0193_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0194_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0195_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0196_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0197_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0198_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0199_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0200_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0201_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0202_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0203_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0204_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0205_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0206_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0207_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0208_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0209_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0210_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0211_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0212_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0213_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0214_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0215_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0216_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0217_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0218_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0219_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0220_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0221_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0222_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0223_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0224_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0225_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0226_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0227_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0228_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0229_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0230_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0231_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0232_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0233_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0234_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0235_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0236_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0237_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0238_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0239_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0240_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0241_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0242_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0243_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0244_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0245_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0246_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0247_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0248_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0249_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0250_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0251_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0252_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0253_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0254_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0255_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0256_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0257_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0258_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0259_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0260_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0261_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0262_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0263_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0264_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0265_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0266_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0267_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0268_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0269_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0270_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0271_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0272_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0273_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0274_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0275_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0276_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0277_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0278_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0279_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0280_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0281_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0282_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0283_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0284_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0285_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0286_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0287_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0288_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0289_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0290_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0291_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0292_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0293_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0294_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0295_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0296_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0297_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0298_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0299_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0300_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0301_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0302_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0303_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0304_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0305_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0306_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0307_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0308_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0309_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0310_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0311_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0312_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0313_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0314_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0315_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0316_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0317_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0318_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0319_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0320_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0321_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0322_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0323_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0324_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0325_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0326_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0327_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0328_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0329_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0330_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0331_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0332_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0333_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0334_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0335_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0336_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0337_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0338_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0339_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0340_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0341_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0342_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0343_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0344_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0345_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0346_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0347_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0348_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0349_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0350_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0351_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0352_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0353_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0354_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0355_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0356_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0357_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0358_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0359_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0360_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0361_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0362_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0363_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0364_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0365_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0366_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0367_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0368_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0369_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0370_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0371_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0372_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0373_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0374_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0375_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0376_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0377_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0378_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0379_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0380_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0381_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0382_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0383_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0384_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0385_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0386_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0387_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0388_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0389_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0390_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0391_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0392_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0393_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0394_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0395_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0396_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0397_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0398_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0399_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0400_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0401_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0402_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0403_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0404_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0405_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0406_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0407_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0408_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0409_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0410_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0411_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0412_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0413_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0414_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0415_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0416_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0417_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0418_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0419_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0420_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0421_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0422_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0423_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0424_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0425_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0426_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0427_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0428_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0429_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0430_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0431_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0432_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0433_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0434_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0435_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0436_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0437_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0438_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0439_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0440_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0441_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0442_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0443_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0444_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0445_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0446_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0447_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0448_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0449_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0450_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0451_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0452_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0453_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0454_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0455_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0456_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0457_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0458_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0459_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0460_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0461_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0462_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0463_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0464_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0465_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0466_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0467_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0468_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0469_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0470_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0471_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0472_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0473_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0474_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0475_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0476_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0477_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0478_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0479_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0480_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0481_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0482_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0483_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0484_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0485_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0486_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0487_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0488_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0489_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0490_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0491_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0492_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0493_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0494_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0495_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0496_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0497_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0498_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0499_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0500_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0501_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0502_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0503_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0504_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0505_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0506_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0507_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0508_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0509_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0510_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0511_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0512_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0513_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0514_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0515_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0516_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0517_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0518_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0519_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0520_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0521_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0522_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0523_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0524_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0525_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0526_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0527_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0528_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0529_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0530_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0531_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0532_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0533_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0534_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0535_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0536_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0537_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0538_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0539_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0540_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0541_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0542_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0543_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0544_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0545_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0546_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0547_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0548_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0549_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0550_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0551_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0552_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0553_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0554_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0555_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0556_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0557_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0558_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0559_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0560_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0561_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0562_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0563_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0564_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0565_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0566_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0567_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0568_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0569_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0570_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0571_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0572_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0573_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0574_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0575_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0576_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0577_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0578_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0579_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0580_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0581_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0582_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0583_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0584_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0585_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0586_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0587_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0588_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0589_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0590_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0591_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0592_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0593_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0594_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0595_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0596_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0597_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0598_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0599_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0600_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0601_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0602_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0603_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0604_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0605_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0606_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0607_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0608_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0609_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0610_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0611_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0612_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0613_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0614_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0615_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0616_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0617_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0618_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0619_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0620_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0621_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0622_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0623_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0624_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0625_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0626_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0627_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0628_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0629_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0630_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0631_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0632_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0633_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0634_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0635_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0636_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0637_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0638_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0639_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0640_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0641_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0642_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0643_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0644_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0645_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0646_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0647_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0648_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0649_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0650_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0651_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0652_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0653_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0654_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0655_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0656_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0657_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0658_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0659_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0660_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0661_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0662_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0663_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0664_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0665_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0666_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0667_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0668_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0669_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0670_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0671_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0672_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0673_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0674_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0675_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0676_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0677_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0678_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0679_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0680_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0681_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0682_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0683_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0684_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0685_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0686_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0687_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0688_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0689_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0690_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0691_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0692_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0693_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0694_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0695_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0696_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0697_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0698_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0699_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0700_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0701_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0702_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0703_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0704_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0705_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0706_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0707_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0708_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0709_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0710_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0711_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0712_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0713_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0714_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0715_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0716_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0717_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0718_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0719_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0720_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0721_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0722_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0723_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0724_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0725_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0726_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0727_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0728_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0729_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0730_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0731_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0732_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0733_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0734_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0735_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0736_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0737_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0738_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0739_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0740_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0741_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0742_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0743_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0744_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0745_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0746_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0747_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0748_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0749_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0750_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0751_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0752_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0753_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0754_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0755_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0756_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0757_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0758_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0759_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0760_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0761_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0762_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0763_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0764_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0765_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0766_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0767_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0768_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0769_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0770_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0771_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0772_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0773_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0774_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0775_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0776_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0777_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0778_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0779_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0780_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0781_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0782_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0783_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0784_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0785_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0786_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0787_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0788_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0789_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0790_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0791_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0792_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0793_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0794_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0795_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0796_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0797_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0798_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0799_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0800_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0801_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0802_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0803_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0804_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0805_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0806_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0807_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0808_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0809_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0810_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0811_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0812_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0813_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0814_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0815_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0816_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0817_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0818_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0819_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0820_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0821_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0822_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0823_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0824_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0825_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0826_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0827_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0828_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0829_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0830_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0831_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0832_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0833_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0834_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0835_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0836_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0837_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0838_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0839_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0840_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0841_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0842_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0843_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0844_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0845_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0846_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0847_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0848_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0849_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0850_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0851_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0852_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0853_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0854_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0855_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0856_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0857_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0858_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0859_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0860_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0861_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0862_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0863_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0864_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0865_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0866_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0867_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0868_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0869_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0870_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0871_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0872_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0873_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0874_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0875_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0876_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0877_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0878_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0879_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0880_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0881_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0882_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0883_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0884_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0885_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0886_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0887_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0888_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0889_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0890_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0891_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0892_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0893_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0894_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0895_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0896_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0897_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0898_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0899_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0900_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0901_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0902_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0903_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0904_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0905_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0906_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0907_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0908_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0909_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0910_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0911_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0912_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0913_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0914_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0915_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0916_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0917_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0918_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0919_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0920_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0921_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0922_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0923_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0924_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0925_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0926_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0927_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0928_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0929_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0930_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0931_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0932_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0933_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0934_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0935_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0936_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0937_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0938_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0939_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0940_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0941_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0942_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0943_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0944_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0945_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0946_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0947_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0948_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0949_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0950_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0951_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0952_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0953_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0954_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0955_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0956_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0957_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0958_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0959_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0960_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0961_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0962_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0963_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0964_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0965_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0966_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0967_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0968_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0969_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0970_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0971_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0972_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [27:0] _0973_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0974_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [13:0] _0975_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [111:0] _0976_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0977_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0978_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0979_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire _0980_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0981_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [111:0] _0982_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0983_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0984_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [111:0] _0985_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0986_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0987_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [111:0] _0988_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0989_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0990_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [111:0] _0991_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0992_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0993_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [111:0] _0994_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0995_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0996_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [111:0] _0997_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0998_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _0999_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [111:0] _1000_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _1001_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3568" *)
  wire [3:0] _1002_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1769" *)
  wire [2:0] _1003_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2132" *)
  wire [2:0] _1004_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1536" *)
  wire [2:0] _1005_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1505" *)
  wire [2:0] _1006_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1240" *)
  wire [3:0] _1007_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1148" *)
  wire [1:0] _1008_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2102" *)
  wire [1:0] _1009_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2151" *)
  wire _1010_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2072" *)
  wire _1011_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5519" *)
  wire _1012_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5641" *)
  wire _1013_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5269" *)
  wire _1014_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2462" *)
  wire [111:0] _1015_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3656" *)
  wire [111:0] _1016_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5086" *)
  wire _1017_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4495" *)
  wire [5:0] _1018_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4410" *)
  wire [115:0] _1019_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4410" *)
  wire [115:0] _1020_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4410" *)
  wire [115:0] _1021_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4410" *)
  wire [115:0] _1022_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4410" *)
  wire [115:0] _1023_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4410" *)
  wire [115:0] _1024_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4410" *)
  wire [115:0] _1025_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4410" *)
  wire [115:0] _1026_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4434" *)
  wire [7:0] _1027_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3961" *)
  wire _1028_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3900" *)
  wire _1029_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2176" *)
  wire [2:0] _1030_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2162" *)
  wire _1031_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2118" *)
  wire [12:0] _1032_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3633" *)
  wire [114:0] _1033_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3610" *)
  wire [114:0] _1034_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3633" *)
  wire [114:0] _1035_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3610" *)
  wire [114:0] _1036_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3633" *)
  wire [114:0] _1037_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3610" *)
  wire [114:0] _1038_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3633" *)
  wire [114:0] _1039_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3610" *)
  wire [114:0] _1040_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3633" *)
  wire [114:0] _1041_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3610" *)
  wire [114:0] _1042_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3633" *)
  wire [114:0] _1043_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3610" *)
  wire [114:0] _1044_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3633" *)
  wire [114:0] _1045_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3610" *)
  wire [114:0] _1046_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3633" *)
  wire [114:0] _1047_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3610" *)
  wire [114:0] _1048_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3778" *)
  wire [5:0] _1049_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4144" *)
  wire [5:0] _1050_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3396" *)
  wire _1051_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3396" *)
  wire _1052_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5028" *)
  wire _1053_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3396" *)
  wire _1054_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5028" *)
  wire _1055_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3396" *)
  wire _1056_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5028" *)
  wire _1057_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4083" *)
  wire [7:0] _1058_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4022" *)
  wire [7:0] _1059_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4268" *)
  wire [7:0] _1060_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4207" *)
  wire [7:0] _1061_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5391" *)
  wire [7:0] _1062_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5147" *)
  wire [7:0] _1063_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1505" *)
  wire _1064_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2272" *)
  wire [2:0] _1065_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2261" *)
  wire _1066_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5580" *)
  wire _1067_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5702" *)
  wire _1068_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5330" *)
  wire _1069_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1859" *)
  wire [2:0] _1070_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1859" *)
  wire [2:0] _1071_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1859" *)
  wire [2:0] _1072_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1859" *)
  wire [2:0] _1073_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1859" *)
  wire [2:0] _1074_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1859" *)
  wire [2:0] _1075_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1859" *)
  wire [2:0] _1076_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6318" *)
  wire [27:0] _1077_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6318" *)
  wire [27:0] _1078_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6318" *)
  wire [27:0] _1079_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6318" *)
  wire [27:0] _1080_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6988" *)
  wire [21:0] _1081_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6988" *)
  wire [21:0] _1082_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6988" *)
  wire [21:0] _1083_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6988" *)
  wire [21:0] _1084_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7642" *)
  wire [15:0] _1085_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7642" *)
  wire [15:0] _1086_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7642" *)
  wire [15:0] _1087_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7642" *)
  wire [15:0] _1088_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5911" *)
  wire _1089_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5985" *)
  wire _1090_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6120" *)
  wire _1091_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6198" *)
  wire [27:0] _1092_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6198" *)
  wire [27:0] _1093_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6198" *)
  wire [27:0] _1094_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6198" *)
  wire [27:0] _1095_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6198" *)
  wire [2:0] _1096_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2094" *)
  wire [12:0] _1097_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5830" *)
  wire [2:0] _1098_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5806" *)
  wire [5:0] _1099_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5922" *)
  wire _1100_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5996" *)
  wire _1101_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6059" *)
  wire _1102_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5848" *)
  wire _1103_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5818" *)
  wire [2:0] _1104_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1384" *)
  wire [2:0] _1105_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1321" *)
  wire [3:0] _1106_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3428" *)
  wire [5:0] _1107_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2051" *)
  wire _1108_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1191" *)
  wire [10:0] _1109_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2061" *)
  wire _1110_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2307" *)
  wire [2:0] _1111_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5028" *)
  wire [2:0] _1112_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5452" *)
  wire [2:0] _1113_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5208" *)
  wire [2:0] _1114_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2292" *)
  wire [2:0] _1115_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2335" *)
  wire _1116_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2351" *)
  wire _1117_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2367" *)
  wire _1118_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2383" *)
  wire _1119_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2399" *)
  wire _1120_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2415" *)
  wire _1121_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2431" *)
  wire _1122_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2447" *)
  wire _1123_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3270" *)
  wire _1124_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3277" *)
  wire _1125_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3284" *)
  wire _1126_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3291" *)
  wire _1127_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3298" *)
  wire _1128_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3305" *)
  wire _1129_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3312" *)
  wire _1130_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3319" *)
  wire _1131_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2648" *)
  wire [2:0] _1132_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2772" *)
  wire [2:0] _1133_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2658" *)
  wire [2:0] _1134_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2833" *)
  wire [2:0] _1135_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2668" *)
  wire [2:0] _1136_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2894" *)
  wire [2:0] _1137_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2678" *)
  wire [2:0] _1138_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2955" *)
  wire [2:0] _1139_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2688" *)
  wire [2:0] _1140_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3016" *)
  wire [2:0] _1141_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2698" *)
  wire [2:0] _1142_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3077" *)
  wire [2:0] _1143_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2708" *)
  wire [2:0] _1144_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3138" *)
  wire [2:0] _1145_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2718" *)
  wire [2:0] _1146_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3199" *)
  wire [2:0] _1147_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1933" *)
  wire _1148_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1933" *)
  wire [1:0] _1149_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1933" *)
  wire [1:0] _1150_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1933" *)
  wire [2:0] _1151_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1933" *)
  wire [2:0] _1152_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4336" *)
  wire _1153_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4352" *)
  wire _1154_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4365" *)
  wire _1155_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1158" *)
  wire [12:0] _1156_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3717" *)
  wire _1157_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2523" *)
  wire _1158_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1203" *)
  wire [7:0] _1159_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3416" *)
  wire [2:0] _1160_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1170" *)
  wire [12:0] _1161_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3839" *)
  wire _1162_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2584" *)
  wire _1163_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1481" *)
  wire [2:0] _1164_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1412" *)
  wire [2:0] _1165_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2241" *)
  wire _1166_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1551" *)
  wire [2:0] _1167_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1551" *)
  wire [2:0] _1168_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1169_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1170_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1171_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1172_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1173_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1174_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1175_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1666" *)
  wire [2:0] _1176_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1666" *)
  wire [2:0] _1177_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1666" *)
  wire [2:0] _1178_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1666" *)
  wire [2:0] _1179_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1666" *)
  wire [2:0] _1180_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1705" *)
  wire [2:0] _1181_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1705" *)
  wire [2:0] _1182_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1705" *)
  wire [2:0] _1183_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1705" *)
  wire [2:0] _1184_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1705" *)
  wire [2:0] _1185_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1705" *)
  wire [2:0] _1186_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1456" *)
  wire [2:0] _1187_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1305" *)
  wire [3:0] _1188_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1412" *)
  wire [2:0] _1189_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2241" *)
  wire _1190_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1551" *)
  wire [2:0] _1191_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1551" *)
  wire [2:0] _1192_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1193_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1194_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1195_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1196_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1197_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1198_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1199_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1666" *)
  wire [2:0] _1200_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1666" *)
  wire [2:0] _1201_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1666" *)
  wire [2:0] _1202_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1666" *)
  wire [2:0] _1203_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1666" *)
  wire [2:0] _1204_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1456" *)
  wire [2:0] _1205_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1305" *)
  wire [3:0] _1206_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1412" *)
  wire [2:0] _1207_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1551" *)
  wire [2:0] _1208_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1551" *)
  wire [2:0] _1209_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1210_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1211_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1212_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1213_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1214_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1215_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1626" *)
  wire [2:0] _1216_;
  wire [1:0] _1217_;
  wire [1:0] _1218_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1551" *)
  wire [2:0] _1219_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1551" *)
  wire [2:0] _1220_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1221_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1222_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1587" *)
  wire [2:0] _1223_;
  wire [1:0] _1224_;
  wire [1:0] _1225_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1551" *)
  wire [2:0] _1226_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1551" *)
  wire [2:0] _1227_;
  wire _1228_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1412" *)
  wire [2:0] _1229_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1153" *)
  wire [1:0] _1230_;
  wire [12:0] _1231_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1177" *)
  wire [12:0] _1232_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1198" *)
  (* unused_bits = "11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _1233_;
  wire [7:0] _1234_;
  wire [3:0] _1235_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1394" *)
  (* unused_bits = "3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _1236_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1522" *)
  wire [2:0] _1237_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1522" *)
  wire [2:0] _1238_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1879" *)
  wire [2:0] _1239_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1888" *)
  wire [2:0] _1240_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1897" *)
  wire [2:0] _1241_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1906" *)
  wire [2:0] _1242_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1915" *)
  wire [2:0] _1243_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1924" *)
  wire [2:0] _1244_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2111" *)
  wire [1:0] _1245_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2126" *)
  wire [12:0] _1246_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2140" *)
  wire [2:0] _1247_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2185" *)
  wire [2:0] _1248_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2280" *)
  wire [2:0] _1249_;
  wire [2:0] _1250_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2655" *)
  wire [2:0] _1251_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2665" *)
  wire [2:0] _1252_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2675" *)
  wire [2:0] _1253_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2685" *)
  wire [2:0] _1254_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2695" *)
  wire [2:0] _1255_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2705" *)
  wire [2:0] _1256_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2715" *)
  wire [2:0] _1257_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2725" *)
  wire [2:0] _1258_;
  wire [2:0] _1259_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3436" *)
  wire [5:0] _1260_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5045" *)
  wire [2:0] _1261_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5813" *)
  wire [5:0] _1262_;
  wire [2:0] _1263_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5838" *)
  (* unused_bits = "3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _1264_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6386" *)
  wire [18:0] _1265_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6387" *)
  wire [18:0] _1266_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6388" *)
  wire [18:0] _1267_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6389" *)
  wire [18:0] _1268_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6611" *)
  wire [10:0] _1269_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6612" *)
  wire [10:0] _1270_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6613" *)
  wire [10:0] _1271_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6614" *)
  wire [10:0] _1272_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6615" *)
  wire [10:0] _1273_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6616" *)
  wire [10:0] _1274_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6617" *)
  wire [10:0] _1275_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6618" *)
  wire [10:0] _1276_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7041" *)
  wire [15:0] _1277_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7042" *)
  wire [15:0] _1278_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7043" *)
  wire [15:0] _1279_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7044" *)
  wire [15:0] _1280_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7266" *)
  wire [7:0] _1281_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7267" *)
  wire [7:0] _1282_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7268" *)
  wire [7:0] _1283_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7269" *)
  wire [7:0] _1284_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7270" *)
  wire [7:0] _1285_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7271" *)
  wire [7:0] _1286_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7272" *)
  wire [7:0] _1287_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7273" *)
  wire [7:0] _1288_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2055" *)
  wire _1289_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2055" *)
  wire _1290_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2065" *)
  wire _1291_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2065" *)
  wire _1292_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2076" *)
  wire _1293_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2076" *)
  wire _1294_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2078" *)
  wire _1295_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2078" *)
  wire _1296_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *)
  wire _1297_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *)
  wire _1298_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *)
  wire _1299_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *)
  wire _1300_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *)
  wire _1301_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *)
  wire _1302_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2182" *)
  wire _1303_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2182" *)
  wire _1304_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2237" *)
  wire _1305_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2265" *)
  wire _1306_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2332" *)
  wire _1307_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2334" *)
  wire _1308_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2348" *)
  wire _1309_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2348" *)
  wire _1310_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2350" *)
  wire _1311_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2364" *)
  wire _1312_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2364" *)
  wire _1313_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2366" *)
  wire _1314_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2380" *)
  wire _1315_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2380" *)
  wire _1316_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2382" *)
  wire _1317_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2396" *)
  wire _1318_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2396" *)
  wire _1319_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2398" *)
  wire _1320_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2412" *)
  wire _1321_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2412" *)
  wire _1322_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2414" *)
  wire _1323_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2428" *)
  wire _1324_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2428" *)
  wire _1325_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2430" *)
  wire _1326_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2444" *)
  wire _1327_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2444" *)
  wire _1328_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2446" *)
  wire _1329_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2654" *)
  wire _1330_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2664" *)
  wire _1331_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2674" *)
  wire _1332_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2684" *)
  wire _1333_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2694" *)
  wire _1334_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2704" *)
  wire _1335_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2714" *)
  wire _1336_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2724" *)
  wire _1337_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3327" *)
  wire _1338_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3327" *)
  wire _1339_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3328" *)
  wire _1340_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3329" *)
  wire _1341_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3330" *)
  wire _1342_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3331" *)
  wire _1343_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3332" *)
  wire _1344_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3333" *)
  wire _1345_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3334" *)
  wire _1346_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3350" *)
  wire _1347_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3350" *)
  wire _1348_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3351" *)
  wire _1349_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3352" *)
  wire _1350_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3353" *)
  wire _1351_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3367" *)
  wire _1352_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3367" *)
  wire _1353_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3368" *)
  wire _1354_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3369" *)
  wire _1355_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3369" *)
  wire _1356_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3370" *)
  wire _1357_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3384" *)
  wire _1358_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3384" *)
  wire _1359_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3385" *)
  wire _1360_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3385" *)
  wire _1361_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3386" *)
  wire _1362_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3386" *)
  wire _1363_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3387" *)
  wire _1364_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3387" *)
  wire _1365_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3435" *)
  wire _1366_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1367_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1368_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1369_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1370_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1371_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1372_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1373_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1374_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1375_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1376_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1377_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1378_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1379_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1380_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1381_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1382_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1383_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1384_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1385_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1386_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1387_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1388_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1389_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1390_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1391_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1392_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1393_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1394_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1395_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1396_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1397_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *)
  wire _1398_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1399_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1400_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1401_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1402_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1403_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1404_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1405_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1406_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1407_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1408_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1409_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1410_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1411_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1412_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1413_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1414_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1415_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1416_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1417_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1418_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1419_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1420_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1421_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1422_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1423_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1424_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1425_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1426_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1427_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1428_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1429_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *)
  wire _1430_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1431_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1432_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1433_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1434_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1435_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1436_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1437_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1438_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1439_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1440_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1441_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1442_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1443_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1444_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1445_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1446_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1447_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1448_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1449_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1450_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1451_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1452_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1453_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1454_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1455_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1456_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1457_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1458_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1459_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1460_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1461_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *)
  wire _1462_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1463_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1464_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1465_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1466_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1467_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1468_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1469_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1470_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1471_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1472_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1473_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1474_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1475_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1476_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1477_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1478_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1479_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1480_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1481_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1482_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1483_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1484_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1485_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1486_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1487_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1488_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1489_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1490_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1491_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1492_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1493_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _1494_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1495_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1496_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1497_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1498_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1499_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1500_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1501_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1502_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1503_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1504_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1505_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1506_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1507_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1508_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1509_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1510_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1511_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1512_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1513_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1514_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1515_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1516_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1517_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1518_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1519_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1520_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1521_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1522_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1523_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1524_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1525_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire _1526_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1527_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1528_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1529_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1530_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1531_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1532_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1533_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1534_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1535_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1536_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1537_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1538_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1539_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1540_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1541_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1542_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1543_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1544_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1545_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1546_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1547_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1548_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1549_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1550_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1551_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1552_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1553_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1554_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1555_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1556_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1557_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire _1558_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1559_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1560_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1561_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1562_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1563_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1564_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1565_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1566_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1567_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1568_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1569_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1570_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1571_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1572_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1573_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1574_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1575_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1576_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1577_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1578_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1579_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1580_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1581_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1582_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1583_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1584_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1585_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1586_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1587_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1588_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1589_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *)
  wire _1590_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1591_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1592_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1593_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1594_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1595_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1596_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1597_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1598_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1599_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1600_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1601_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1602_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1603_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1604_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1605_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1606_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1607_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1608_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1609_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1610_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1611_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1612_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1613_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1614_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1615_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1616_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1617_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1618_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1619_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1620_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1621_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *)
  wire _1622_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1623_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1624_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1625_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1626_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1627_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1628_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1629_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1630_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1631_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1632_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1633_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1634_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1635_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1636_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1637_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1638_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1639_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1640_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1641_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1642_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1643_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1644_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1645_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1646_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1647_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1648_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1649_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1650_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1651_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1652_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1653_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *)
  wire _1654_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *)
  wire _1655_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *)
  wire _1656_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *)
  wire _1657_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *)
  wire _1658_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *)
  wire _1659_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *)
  wire _1660_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *)
  wire _1661_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *)
  wire _1662_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *)
  wire _1663_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *)
  wire _1664_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *)
  wire _1665_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *)
  wire _1666_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *)
  wire _1667_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *)
  wire _1668_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *)
  wire _1669_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *)
  wire _1670_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _1671_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _1672_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _1673_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _1674_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _1675_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _1676_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _1677_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _1678_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _1679_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _1680_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _1681_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _1682_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _1683_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _1684_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _1685_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _1686_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _1687_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _1688_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _1689_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _1690_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _1691_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _1692_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _1693_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _1694_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _1695_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _1696_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _1697_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _1698_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _1699_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _1700_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _1701_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _1702_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3621" *)
  wire _1703_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4148" *)
  wire _1704_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4351" *)
  wire _1705_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4364" *)
  wire _1706_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4370" *)
  wire _1707_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4377" *)
  wire _1708_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4566" *)
  wire [7:0] _1709_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5041" *)
  wire _1710_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5041" *)
  wire _1711_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5041" *)
  wire _1712_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5061" *)
  wire _1713_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5062" *)
  wire _1714_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5063" *)
  wire _1715_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5064" *)
  wire _1716_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5065" *)
  wire _1717_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5066" *)
  wire _1718_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5067" *)
  wire _1719_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5068" *)
  wire _1720_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5073" *)
  wire _1721_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5074" *)
  wire _1722_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5075" *)
  wire _1723_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5076" *)
  wire _1724_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5081" *)
  wire _1725_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5082" *)
  wire _1726_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5083" *)
  wire _1727_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5084" *)
  wire _1728_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5090" *)
  wire _1729_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5395" *)
  wire _1730_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5456" *)
  wire _1731_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5764" *)
  wire _1732_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5764" *)
  wire _1733_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5764" *)
  wire _1734_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5765" *)
  wire _1735_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5765" *)
  wire _1736_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5766" *)
  wire _1737_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5766" *)
  wire _1738_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5767" *)
  wire _1739_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5767" *)
  wire _1740_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5768" *)
  wire _1741_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5768" *)
  wire _1742_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5769" *)
  wire _1743_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5769" *)
  wire _1744_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5770" *)
  wire _1745_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5770" *)
  wire _1746_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5771" *)
  wire _1747_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5771" *)
  wire _1748_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5775" *)
  wire _1749_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5776" *)
  wire _1750_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5777" *)
  wire _1751_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5778" *)
  wire _1752_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5779" *)
  wire _1753_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5780" *)
  wire _1754_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5783" *)
  wire _1755_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5784" *)
  wire _1756_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5785" *)
  wire _1757_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5786" *)
  wire _1758_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5787" *)
  wire _1759_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5788" *)
  wire _1760_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5789" *)
  wire _1761_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5791" *)
  wire [114:0] _1762_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5792" *)
  wire [114:0] _1763_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5793" *)
  wire [114:0] _1764_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5794" *)
  wire [114:0] _1765_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5795" *)
  wire [114:0] _1766_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5796" *)
  wire [114:0] _1767_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5797" *)
  wire [114:0] _1768_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5798" *)
  wire [114:0] _1769_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5816" *)
  wire _1770_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5828" *)
  wire _1771_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5835" *)
  wire _1772_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5837" *)
  wire _1773_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5841" *)
  wire _1774_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5845" *)
  wire _1775_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6132" *)
  wire [7:0] _1776_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6132" *)
  wire [7:0] _1777_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6134" *)
  wire _1778_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6134" *)
  wire _1779_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6134" *)
  wire _1780_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6135" *)
  wire _1781_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6135" *)
  wire _1782_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6135" *)
  wire _1783_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6136" *)
  wire _1784_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6136" *)
  wire _1785_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6136" *)
  wire _1786_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6137" *)
  wire _1787_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6137" *)
  wire _1788_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6137" *)
  wire _1789_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6138" *)
  wire _1790_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6138" *)
  wire _1791_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6138" *)
  wire _1792_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6139" *)
  wire _1793_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6139" *)
  wire _1794_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6139" *)
  wire _1795_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6140" *)
  wire _1796_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6140" *)
  wire _1797_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6140" *)
  wire _1798_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6141" *)
  wire _1799_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6141" *)
  wire _1800_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6141" *)
  wire _1801_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6145" *)
  wire _1802_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6145" *)
  wire _1803_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6146" *)
  wire _1804_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6146" *)
  wire _1805_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6147" *)
  wire _1806_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6147" *)
  wire _1807_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6148" *)
  wire _1808_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6148" *)
  wire _1809_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6149" *)
  wire _1810_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6149" *)
  wire _1811_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6150" *)
  wire _1812_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6150" *)
  wire _1813_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6153" *)
  wire _1814_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6153" *)
  wire _1815_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6154" *)
  wire _1816_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6154" *)
  wire _1817_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6155" *)
  wire _1818_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6155" *)
  wire _1819_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6156" *)
  wire _1820_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6156" *)
  wire _1821_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6157" *)
  wire _1822_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6157" *)
  wire _1823_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6158" *)
  wire _1824_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6158" *)
  wire _1825_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6159" *)
  wire _1826_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6159" *)
  wire _1827_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6325" *)
  wire _1828_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6374" *)
  wire _1829_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6375" *)
  wire _1830_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6376" *)
  wire _1831_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6377" *)
  wire _1832_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6378" *)
  wire _1833_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6379" *)
  wire _1834_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6380" *)
  wire _1835_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6381" *)
  wire _1836_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6587" *)
  wire _1837_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6588" *)
  wire _1838_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6589" *)
  wire _1839_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6590" *)
  wire _1840_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6591" *)
  wire _1841_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6592" *)
  wire _1842_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6593" *)
  wire _1843_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6594" *)
  wire _1844_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6595" *)
  wire _1845_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6596" *)
  wire _1846_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6597" *)
  wire _1847_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6598" *)
  wire _1848_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6599" *)
  wire _1849_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6600" *)
  wire _1850_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6601" *)
  wire _1851_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6602" *)
  wire _1852_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7029" *)
  wire _1853_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7030" *)
  wire _1854_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7031" *)
  wire _1855_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7032" *)
  wire _1856_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7033" *)
  wire _1857_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7034" *)
  wire _1858_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7035" *)
  wire _1859_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7036" *)
  wire _1860_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7242" *)
  wire _1861_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7243" *)
  wire _1862_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7244" *)
  wire _1863_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7245" *)
  wire _1864_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7246" *)
  wire _1865_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7247" *)
  wire _1866_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7248" *)
  wire _1867_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7249" *)
  wire _1868_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7250" *)
  wire _1869_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7251" *)
  wire _1870_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7252" *)
  wire _1871_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7253" *)
  wire _1872_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7254" *)
  wire _1873_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7255" *)
  wire _1874_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7256" *)
  wire _1875_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7257" *)
  wire _1876_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7784" *)
  wire _1877_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7785" *)
  wire _1878_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7786" *)
  wire _1879_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7787" *)
  wire _1880_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7788" *)
  wire _1881_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7789" *)
  wire _1882_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7790" *)
  wire _1883_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7791" *)
  wire _1884_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7953" *)
  wire _1885_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7954" *)
  wire _1886_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7955" *)
  wire _1887_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7956" *)
  wire _1888_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7957" *)
  wire _1889_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7958" *)
  wire _1890_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7959" *)
  wire _1891_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7960" *)
  wire _1892_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7963" *)
  wire _1893_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7963" *)
  wire _1894_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8023" *)
  wire [114:0] _1895_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8024" *)
  wire [114:0] _1896_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8025" *)
  wire [114:0] _1897_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8026" *)
  wire [114:0] _1898_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8027" *)
  wire [114:0] _1899_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8028" *)
  wire [114:0] _1900_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8029" *)
  wire [114:0] _1901_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8030" *)
  wire [114:0] _1902_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8031" *)
  wire [114:0] _1903_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8032" *)
  wire [114:0] _1904_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8033" *)
  wire [114:0] _1905_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8034" *)
  wire [114:0] _1906_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8035" *)
  wire [114:0] _1907_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8036" *)
  wire [114:0] _1908_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8037" *)
  wire [114:0] _1909_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8038" *)
  wire [114:0] _1910_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8788" *)
  wire _1911_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8789" *)
  wire _1912_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1299" *)
  (* unused_bits = "3 4 5 6 7" *)
  wire [8:0] _1913_;
  wire [2:0] _1914_;
  wire [2:0] _1915_;
  wire [2:0] _1916_;
  wire [2:0] _1917_;
  wire [2:0] _1918_;
  wire [2:0] _1919_;
  wire [2:0] _1920_;
  wire [2:0] _1921_;
  wire [2:0] _1922_;
  wire [2:0] _1923_;
  wire [2:0] _1924_;
  wire [2:0] _1925_;
  wire [2:0] _1926_;
  wire [2:0] _1927_;
  wire [2:0] _1928_;
  wire [2:0] _1929_;
  wire [2:0] _1930_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1504" *)
  (* unused_bits = "4" *)
  wire [4:0] _1931_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [31:0] _1932_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [31:0] _1933_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [31:0] _1934_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [31:0] _1935_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [31:0] _1936_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [31:0] _1937_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [31:0] _1938_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [31:0] _1939_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _1940_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _1941_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _1942_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _1943_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _1944_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _1945_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _1946_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _1947_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [31:0] _1948_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [31:0] _1949_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [31:0] _1950_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [31:0] _1951_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [31:0] _1952_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [31:0] _1953_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [31:0] _1954_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [31:0] _1955_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _1956_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _1957_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _1958_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _1959_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _1960_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _1961_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _1962_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _1963_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _1964_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [31:0] _1965_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [31:0] _1966_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [31:0] _1967_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [31:0] _1968_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [31:0] _1969_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [31:0] _1970_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [31:0] _1971_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [31:0] _1972_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _1973_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _1974_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _1975_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _1976_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _1977_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _1978_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _1979_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _1980_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [31:0] _1981_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [31:0] _1982_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [31:0] _1983_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [31:0] _1984_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [31:0] _1985_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [31:0] _1986_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [31:0] _1987_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [31:0] _1988_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _1989_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _1990_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _1991_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _1992_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _1993_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _1994_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _1995_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _1996_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _1997_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _1998_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _1999_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _2000_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _2001_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _2002_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _2003_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _2004_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _2005_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _2006_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _2007_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _2008_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _2009_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _2010_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1168" *)
  wire _2011_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1201" *)
  wire _2012_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1213" *)
  wire _2013_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1218" *)
  wire _2014_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1302" *)
  wire _2015_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1325" *)
  wire _2016_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1465" *)
  wire _2017_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1467" *)
  wire _2018_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1469" *)
  wire _2019_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1471" *)
  wire _2020_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1473" *)
  wire _2021_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1486" *)
  wire _2022_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1562" *)
  wire _2023_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1563" *)
  wire _2024_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1566" *)
  wire _2025_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1569" *)
  wire _2026_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1572" *)
  wire _2027_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1575" *)
  wire _2028_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1598" *)
  wire _2029_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1637" *)
  wire _2030_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1677" *)
  wire _2031_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1716" *)
  wire _2032_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1751" *)
  wire _2033_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *)
  wire _2034_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *)
  wire _2035_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *)
  wire _2036_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *)
  wire _2037_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *)
  wire _2038_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *)
  wire _2039_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *)
  wire _2040_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *)
  wire _2041_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *)
  wire _2042_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *)
  wire _2043_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *)
  wire _2044_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *)
  wire _2045_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *)
  wire _2046_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *)
  wire _2047_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *)
  wire _2048_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *)
  wire _2049_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *)
  wire _2050_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *)
  wire _2051_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *)
  wire _2052_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *)
  wire _2053_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *)
  wire _2054_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *)
  wire _2055_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *)
  wire _2056_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *)
  wire _2057_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *)
  wire _2058_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *)
  wire _2059_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *)
  wire _2060_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *)
  wire _2061_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *)
  wire _2062_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *)
  wire _2063_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *)
  wire _2064_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *)
  wire _2065_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *)
  wire _2066_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *)
  wire _2067_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *)
  wire _2068_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *)
  wire _2069_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *)
  wire _2070_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *)
  wire _2071_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *)
  wire _2072_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *)
  wire _2073_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *)
  wire _2074_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *)
  wire _2075_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *)
  wire _2076_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *)
  wire _2077_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *)
  wire _2078_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *)
  wire _2079_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *)
  wire _2080_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *)
  wire _2081_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *)
  wire _2082_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *)
  wire _2083_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *)
  wire _2084_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *)
  wire _2085_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *)
  wire _2086_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *)
  wire _2087_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *)
  wire _2088_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *)
  wire _2089_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *)
  wire _2090_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *)
  wire _2091_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *)
  wire _2092_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *)
  wire _2093_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *)
  wire _2094_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *)
  wire _2095_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *)
  wire _2096_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *)
  wire _2097_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *)
  wire _2098_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *)
  wire _2099_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *)
  wire _2100_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *)
  wire _2101_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *)
  wire _2102_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *)
  wire _2103_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *)
  wire _2104_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *)
  wire _2105_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *)
  wire _2106_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *)
  wire _2107_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *)
  wire _2108_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *)
  wire _2109_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *)
  wire _2110_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *)
  wire _2111_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *)
  wire _2112_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *)
  wire _2113_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *)
  wire _2114_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *)
  wire _2115_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *)
  wire _2116_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *)
  wire _2117_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *)
  wire _2118_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *)
  wire _2119_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *)
  wire _2120_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *)
  wire _2121_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *)
  wire _2122_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *)
  wire _2123_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *)
  wire _2124_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *)
  wire _2125_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *)
  wire _2126_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *)
  wire _2127_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *)
  wire _2128_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *)
  wire _2129_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *)
  wire _2130_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *)
  wire _2131_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *)
  wire _2132_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *)
  wire _2133_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *)
  wire _2134_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *)
  wire _2135_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *)
  wire _2136_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *)
  wire _2137_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *)
  wire _2138_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *)
  wire _2139_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *)
  wire _2140_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *)
  wire _2141_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *)
  wire _2142_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *)
  wire _2143_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *)
  wire _2144_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *)
  wire _2145_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *)
  wire _2146_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *)
  wire _2147_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *)
  wire _2148_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *)
  wire _2149_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *)
  wire _2150_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *)
  wire _2151_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *)
  wire _2152_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *)
  wire _2153_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *)
  wire _2154_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *)
  wire _2155_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *)
  wire _2156_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *)
  wire _2157_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *)
  wire _2158_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *)
  wire _2159_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *)
  wire _2160_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *)
  wire _2161_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *)
  wire _2162_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *)
  wire _2163_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *)
  wire _2164_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *)
  wire _2165_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *)
  wire _2166_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *)
  wire _2167_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *)
  wire _2168_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *)
  wire _2169_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *)
  wire _2170_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *)
  wire _2171_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *)
  wire _2172_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *)
  wire _2173_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *)
  wire _2174_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *)
  wire _2175_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *)
  wire _2176_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *)
  wire _2177_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *)
  wire _2178_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *)
  wire _2179_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *)
  wire _2180_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *)
  wire _2181_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *)
  wire _2182_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *)
  wire _2183_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *)
  wire _2184_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *)
  wire _2185_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *)
  wire _2186_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *)
  wire _2187_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *)
  wire _2188_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *)
  wire _2189_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *)
  wire _2190_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *)
  wire _2191_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *)
  wire _2192_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *)
  wire _2193_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *)
  wire _2194_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *)
  wire _2195_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1870" *)
  wire _2196_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1878" *)
  wire _2197_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1886" *)
  wire _2198_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1894" *)
  wire _2199_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1902" *)
  wire _2200_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1910" *)
  wire _2201_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1918" *)
  wire _2202_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1934" *)
  wire _2203_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1940" *)
  wire _2204_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1941" *)
  wire _2205_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1954" *)
  wire _2206_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1961" *)
  wire _2207_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1974" *)
  wire _2208_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1981" *)
  wire _2209_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1994" *)
  wire _2210_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2007" *)
  wire _2211_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2020" *)
  wire _2212_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2033" *)
  wire _2213_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2117" *)
  wire _2214_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2131" *)
  wire _2215_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2145" *)
  wire _2216_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2182" *)
  wire _2217_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2182" *)
  wire _2218_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2252" *)
  wire _2219_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2254" *)
  wire _2220_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2256" *)
  wire _2221_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2258" *)
  wire _2222_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2285" *)
  wire _2223_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2287" *)
  wire _2224_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2334" *)
  wire _2225_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2348" *)
  wire _2226_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2350" *)
  wire _2227_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2364" *)
  wire _2228_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2366" *)
  wire _2229_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2380" *)
  wire _2230_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2382" *)
  wire _2231_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2396" *)
  wire _2232_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2398" *)
  wire _2233_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2412" *)
  wire _2234_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2414" *)
  wire _2235_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2428" *)
  wire _2236_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2430" *)
  wire _2237_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2444" *)
  wire _2238_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2446" *)
  wire _2239_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3327" *)
  wire _2240_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3328" *)
  wire _2241_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3329" *)
  wire _2242_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3330" *)
  wire _2243_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3331" *)
  wire _2244_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3332" *)
  wire _2245_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3333" *)
  wire _2246_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3334" *)
  wire _2247_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3405" *)
  wire _2248_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3405" *)
  wire _2249_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3426" *)
  wire _2250_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3440" *)
  wire _2251_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4148" *)
  wire _2252_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5053" *)
  wire _2253_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5054" *)
  wire _2254_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5055" *)
  wire _2255_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5056" *)
  wire _2256_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5057" *)
  wire _2257_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5058" *)
  wire _2258_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5059" *)
  wire _2259_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5060" *)
  wire _2260_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5090" *)
  wire _2261_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5151" *)
  wire _2262_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5395" *)
  wire _2263_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5456" *)
  wire _2264_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5764" *)
  wire _2265_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5768" *)
  wire _2266_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5777" *)
  wire _2267_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5779" *)
  wire _2268_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5786" *)
  wire _2269_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5787" *)
  wire _2270_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5788" *)
  wire _2271_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5789" *)
  wire _2272_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5816" *)
  wire _2273_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5828" *)
  wire _2274_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5841" *)
  wire _2275_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6134" *)
  wire _2276_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6138" *)
  wire _2277_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6147" *)
  wire _2278_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6149" *)
  wire _2279_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6156" *)
  wire _2280_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6157" *)
  wire _2281_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6158" *)
  wire _2282_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6159" *)
  wire _2283_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1236" *)
  wire _2284_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1279" *)
  wire _2285_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1280" *)
  wire _2286_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1390" *)
  wire _2287_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1520" *)
  wire _2288_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2331" *)
  wire _2289_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2347" *)
  wire _2290_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2363" *)
  wire _2291_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2379" *)
  wire _2292_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2395" *)
  wire _2293_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2411" *)
  wire _2294_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2427" *)
  wire _2295_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2443" *)
  wire _2296_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2258" *)
  wire _2297_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2298_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2299_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2300_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2301_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2302_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2303_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2304_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2305_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2306_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2307_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2308_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2309_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2310_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2311_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2312_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2313_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2314_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2315_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2316_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2317_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2318_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2319_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2320_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2321_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2322_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2323_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2324_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2325_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2326_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2327_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2328_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2329_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1396" *)
  wire _2330_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2098" *)
  wire _2331_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1422" *)
  wire _2332_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1424" *)
  wire _2333_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1426" *)
  wire _2334_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1428" *)
  wire _2335_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1430" *)
  wire _2336_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1432" *)
  wire _2337_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1434" *)
  wire _2338_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1440" *)
  wire _2339_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *)
  wire _2340_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2166" *)
  wire _2341_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6220" *)
  wire _2342_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1139" *)
  wire _2343_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1140" *)
  wire _2344_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1301" *)
  wire _2345_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1440" *)
  wire _2346_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2076" *)
  wire _2347_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *)
  wire _2348_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *)
  wire _2349_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *)
  wire _2350_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2332" *)
  wire _2351_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2348" *)
  wire _2352_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2353_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2354_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2355_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2356_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2357_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2358_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2359_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2360_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2361_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2362_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2363_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2364_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2365_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2366_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2367_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2368_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2369_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2370_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2371_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2372_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2373_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2374_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2375_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2376_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2377_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2378_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2379_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2380_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2381_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2382_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2383_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2384_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2385_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2386_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2387_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire _2388_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2389_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2390_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2391_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2392_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2393_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2394_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2395_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2396_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2397_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2398_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2399_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2400_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2401_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2402_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2403_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2404_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2405_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2406_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2407_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2408_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2409_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2410_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2411_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2412_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2413_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2414_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2415_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2416_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2417_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2418_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2419_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2420_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2421_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4330" *)
  wire _2422_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4347" *)
  wire _2423_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4351" *)
  wire _2424_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4351" *)
  wire _2425_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4364" *)
  wire _2426_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4364" *)
  wire _2427_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4370" *)
  wire _2428_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4377" *)
  wire _2429_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4377" *)
  wire _2430_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5847" *)
  wire _2431_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5910" *)
  wire _2432_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5921" *)
  wire _2433_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5995" *)
  wire _2434_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6325" *)
  wire _2435_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6374" *)
  wire _2436_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6374" *)
  wire _2437_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6375" *)
  wire _2438_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6375" *)
  wire _2439_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6376" *)
  wire _2440_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6376" *)
  wire _2441_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6377" *)
  wire _2442_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6377" *)
  wire _2443_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6587" *)
  wire _2444_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6587" *)
  wire _2445_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6588" *)
  wire _2446_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6588" *)
  wire _2447_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6589" *)
  wire _2448_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6589" *)
  wire _2449_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6590" *)
  wire _2450_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6590" *)
  wire _2451_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6591" *)
  wire _2452_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6591" *)
  wire _2453_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6592" *)
  wire _2454_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6592" *)
  wire _2455_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6593" *)
  wire _2456_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6593" *)
  wire _2457_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6594" *)
  wire _2458_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6594" *)
  wire _2459_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7029" *)
  wire _2460_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7029" *)
  wire _2461_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7030" *)
  wire _2462_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7030" *)
  wire _2463_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7031" *)
  wire _2464_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7031" *)
  wire _2465_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7032" *)
  wire _2466_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7032" *)
  wire _2467_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7242" *)
  wire _2468_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7242" *)
  wire _2469_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7243" *)
  wire _2470_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7243" *)
  wire _2471_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7244" *)
  wire _2472_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7244" *)
  wire _2473_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7245" *)
  wire _2474_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7245" *)
  wire _2475_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7246" *)
  wire _2476_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7246" *)
  wire _2477_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7247" *)
  wire _2478_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7247" *)
  wire _2479_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7248" *)
  wire _2480_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7248" *)
  wire _2481_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7249" *)
  wire _2482_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7249" *)
  wire _2483_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7963" *)
  wire _2484_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7963" *)
  wire _2485_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1325" *)
  wire _2486_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *)
  wire _2487_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *)
  wire _2488_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *)
  wire _2489_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *)
  wire _2490_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *)
  wire _2491_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *)
  wire _2492_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *)
  wire _2493_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *)
  wire _2494_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *)
  wire _2495_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *)
  wire _2496_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *)
  wire _2497_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *)
  wire _2498_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *)
  wire _2499_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *)
  wire _2500_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *)
  wire _2501_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *)
  wire _2502_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *)
  wire _2503_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *)
  wire _2504_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *)
  wire _2505_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *)
  wire _2506_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *)
  wire _2507_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *)
  wire _2508_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *)
  wire _2509_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *)
  wire _2510_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *)
  wire _2511_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *)
  wire _2512_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *)
  wire _2513_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *)
  wire _2514_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *)
  wire _2515_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *)
  wire _2516_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *)
  wire _2517_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *)
  wire _2518_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *)
  wire _2519_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *)
  wire _2520_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *)
  wire _2521_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *)
  wire _2522_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *)
  wire _2523_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *)
  wire _2524_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *)
  wire _2525_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *)
  wire _2526_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *)
  wire _2527_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *)
  wire _2528_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *)
  wire _2529_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *)
  wire _2530_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *)
  wire _2531_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *)
  wire _2532_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *)
  wire _2533_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *)
  wire _2534_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *)
  wire _2535_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *)
  wire _2536_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *)
  wire _2537_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *)
  wire _2538_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *)
  wire _2539_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *)
  wire _2540_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *)
  wire _2541_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *)
  wire _2542_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *)
  wire _2543_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *)
  wire _2544_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *)
  wire _2545_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *)
  wire _2546_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *)
  wire _2547_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *)
  wire _2548_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *)
  wire _2549_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *)
  wire _2550_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *)
  wire _2551_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *)
  wire _2552_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *)
  wire _2553_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *)
  wire _2554_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *)
  wire _2555_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *)
  wire _2556_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *)
  wire _2557_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *)
  wire _2558_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *)
  wire _2559_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *)
  wire _2560_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *)
  wire _2561_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *)
  wire _2562_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *)
  wire _2563_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *)
  wire _2564_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *)
  wire _2565_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *)
  wire _2566_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *)
  wire _2567_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *)
  wire _2568_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *)
  wire _2569_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *)
  wire _2570_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *)
  wire _2571_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *)
  wire _2572_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *)
  wire _2573_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *)
  wire _2574_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *)
  wire _2575_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *)
  wire _2576_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *)
  wire _2577_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *)
  wire _2578_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *)
  wire _2579_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *)
  wire _2580_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *)
  wire _2581_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *)
  wire _2582_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *)
  wire _2583_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *)
  wire _2584_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *)
  wire _2585_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *)
  wire _2586_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *)
  wire _2587_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *)
  wire _2588_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *)
  wire _2589_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *)
  wire _2590_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *)
  wire _2591_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *)
  wire _2592_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *)
  wire _2593_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *)
  wire _2594_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *)
  wire _2595_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *)
  wire _2596_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *)
  wire _2597_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *)
  wire _2598_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *)
  wire _2599_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *)
  wire _2600_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *)
  wire _2601_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *)
  wire _2602_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *)
  wire _2603_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *)
  wire _2604_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *)
  wire _2605_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *)
  wire _2606_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *)
  wire _2607_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *)
  wire _2608_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *)
  wire _2609_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *)
  wire _2610_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *)
  wire _2611_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *)
  wire _2612_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *)
  wire _2613_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *)
  wire _2614_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *)
  wire _2615_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1981" *)
  wire _2616_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2007" *)
  wire _2617_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2033" *)
  wire _2618_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2076" *)
  wire _2619_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2078" *)
  wire _2620_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *)
  wire _2621_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2182" *)
  wire _2622_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2313" *)
  wire _2623_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2764" *)
  wire [2:0] _2624_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2764" *)
  wire [2:0] _2625_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2766" *)
  wire [2:0] _2626_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2768" *)
  wire [2:0] _2627_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2768" *)
  wire [2:0] _2628_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2770" *)
  wire [2:0] _2629_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3412" *)
  wire [7:0] _2630_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3412" *)
  wire [7:0] _2631_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3413" *)
  wire [7:0] _2632_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3413" *)
  wire [7:0] _2633_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3420" *)
  wire _2634_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3420" *)
  wire _2635_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3432" *)
  wire _2636_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3432" *)
  wire _2637_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2638_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2639_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2640_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2641_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2642_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2643_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2644_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire _2645_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2646_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2647_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2648_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2649_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2650_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2651_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2652_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire _2653_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2654_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2655_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2656_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2657_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2658_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2659_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2660_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire _2661_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2662_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2663_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2664_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2665_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2666_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2667_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2668_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire _2669_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4333" *)
  wire _2670_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4582" *)
  wire _2671_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4592" *)
  wire _2672_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4602" *)
  wire _2673_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4612" *)
  wire _2674_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4622" *)
  wire _2675_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4632" *)
  wire _2676_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4642" *)
  wire _2677_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4652" *)
  wire _2678_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5041" *)
  wire _2679_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5052" *)
  wire _2680_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5085" *)
  wire [7:0] _2681_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5764" *)
  wire _2682_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5790" *)
  wire [7:0] _2683_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5792" *)
  wire [114:0] _2684_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5793" *)
  wire [114:0] _2685_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5794" *)
  wire [114:0] _2686_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5795" *)
  wire [114:0] _2687_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5796" *)
  wire [114:0] _2688_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5797" *)
  wire [114:0] _2689_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5810" *)
  wire _2690_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5835" *)
  wire _2691_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5845" *)
  wire _2692_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5847" *)
  wire _2693_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6160" *)
  wire [7:0] _2694_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6160" *)
  wire [7:0] _2695_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6374" *)
  wire _2696_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6375" *)
  wire _2697_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6376" *)
  wire _2698_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6377" *)
  wire _2699_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6587" *)
  wire _2700_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6588" *)
  wire _2701_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6589" *)
  wire _2702_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6590" *)
  wire _2703_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6591" *)
  wire _2704_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6592" *)
  wire _2705_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6593" *)
  wire _2706_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6594" *)
  wire _2707_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7029" *)
  wire _2708_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7030" *)
  wire _2709_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7031" *)
  wire _2710_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7032" *)
  wire _2711_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7242" *)
  wire _2712_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7243" *)
  wire _2713_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7244" *)
  wire _2714_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7245" *)
  wire _2715_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7246" *)
  wire _2716_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7247" *)
  wire _2717_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7248" *)
  wire _2718_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7249" *)
  wire _2719_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8025" *)
  wire [114:0] _2720_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8026" *)
  wire [114:0] _2721_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8027" *)
  wire [114:0] _2722_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8028" *)
  wire [114:0] _2723_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8029" *)
  wire [114:0] _2724_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8030" *)
  wire [114:0] _2725_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8033" *)
  wire [114:0] _2726_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8034" *)
  wire [114:0] _2727_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8035" *)
  wire [114:0] _2728_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8036" *)
  wire [114:0] _2729_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8037" *)
  wire [114:0] _2730_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8038" *)
  wire [114:0] _2731_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8762" *)
  wire [7:0] _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire [15:0] _2740_;
  wire [15:0] _2741_;
  wire [15:0] _2742_;
  wire [15:0] _2743_;
  wire [15:0] _2744_;
  wire [15:0] _2745_;
  wire [15:0] _2746_;
  wire [15:0] _2747_;
  wire [15:0] _2748_;
  wire [15:0] _2749_;
  wire [15:0] _2750_;
  wire [15:0] _2751_;
  wire [21:0] _2752_;
  wire [21:0] _2753_;
  wire [21:0] _2754_;
  wire [21:0] _2755_;
  wire [21:0] _2756_;
  wire [21:0] _2757_;
  wire [21:0] _2758_;
  wire [21:0] _2759_;
  wire [21:0] _2760_;
  wire [21:0] _2761_;
  wire [21:0] _2762_;
  wire [21:0] _2763_;
  wire [27:0] _2764_;
  wire [27:0] _2765_;
  wire [27:0] _2766_;
  wire [27:0] _2767_;
  wire [27:0] _2768_;
  wire [27:0] _2769_;
  wire [27:0] _2770_;
  wire [27:0] _2771_;
  wire [27:0] _2772_;
  wire [27:0] _2773_;
  wire [27:0] _2774_;
  wire [27:0] _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire [2:0] _2794_;
  wire [2:0] _2795_;
  wire [5:0] _2796_;
  wire [2:0] _2797_;
  wire [2:0] _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire [5:0] _2802_;
  wire [2:0] _2803_;
  wire [2:0] _2804_;
  wire [2:0] _2805_;
  wire [2:0] _2806_;
  wire [2:0] _2807_;
  wire [2:0] _2808_;
  wire [2:0] _2809_;
  wire [2:0] _2810_;
  wire [2:0] _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire [2:0] _2828_;
  wire [2:0] _2829_;
  wire [2:0] _2830_;
  wire [2:0] _2831_;
  wire [2:0] _2832_;
  wire [2:0] _2833_;
  wire _2834_;
  wire [2:0] _2835_;
  wire [2:0] _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire [2:0] _2840_;
  wire [2:0] _2841_;
  wire [12:0] _2842_;
  wire [12:0] _2843_;
  wire [1:0] _2844_;
  wire [1:0] _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire [2:0] _2850_;
  wire [2:0] _2851_;
  wire [2:0] _2852_;
  wire [2:0] _2853_;
  wire [2:0] _2854_;
  wire [2:0] _2855_;
  wire [2:0] _2856_;
  wire [2:0] _2857_;
  wire [2:0] _2858_;
  wire [2:0] _2859_;
  wire [2:0] _2860_;
  wire [2:0] _2861_;
  wire [1:0] _2862_;
  wire [1:0] _2863_;
  wire [1:0] _2864_;
  wire [1:0] _2865_;
  wire [1:0] _2866_;
  wire [1:0] _2867_;
  wire [1:0] _2868_;
  wire [1:0] _2869_;
  wire [1:0] _2870_;
  wire [1:0] _2871_;
  wire [1:0] _2872_;
  wire [1:0] _2873_;
  wire [1:0] _2874_;
  wire [1:0] _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire [2:0] _2887_;
  wire [2:0] _2888_;
  wire [2:0] _2889_;
  wire [2:0] _2890_;
  wire [2:0] _2891_;
  wire [2:0] _2892_;
  wire [2:0] _2893_;
  wire [2:0] _2894_;
  wire [2:0] _2895_;
  wire [2:0] _2896_;
  wire [2:0] _2897_;
  wire [2:0] _2898_;
  wire [2:0] _2899_;
  wire [2:0] _2900_;
  wire [2:0] _2901_;
  wire [2:0] _2902_;
  wire [2:0] _2903_;
  wire [2:0] _2904_;
  wire [2:0] _2905_;
  wire [2:0] _2906_;
  wire [2:0] _2907_;
  wire [2:0] _2908_;
  wire [2:0] _2909_;
  wire [2:0] _2910_;
  wire [2:0] _2911_;
  wire [2:0] _2912_;
  wire [2:0] _2913_;
  wire [2:0] _2914_;
  wire [2:0] _2915_;
  wire [2:0] _2916_;
  wire [2:0] _2917_;
  wire [2:0] _2918_;
  wire [2:0] _2919_;
  wire [2:0] _2920_;
  wire [2:0] _2921_;
  wire [2:0] _2922_;
  wire [2:0] _2923_;
  wire [2:0] _2924_;
  wire [2:0] _2925_;
  wire [2:0] _2926_;
  wire [2:0] _2927_;
  wire [2:0] _2928_;
  wire [2:0] _2929_;
  wire [2:0] _2930_;
  wire [2:0] _2931_;
  wire [2:0] _2932_;
  wire [2:0] _2933_;
  wire [2:0] _2934_;
  wire [2:0] _2935_;
  wire [2:0] _2936_;
  wire [2:0] _2937_;
  wire [2:0] _2938_;
  wire [2:0] _2939_;
  wire [2:0] _2940_;
  wire [2:0] _2941_;
  wire [2:0] _2942_;
  wire [2:0] _2943_;
  wire [2:0] _2944_;
  wire [2:0] _2945_;
  wire [2:0] _2946_;
  wire [2:0] _2947_;
  wire [2:0] _2948_;
  wire [2:0] _2949_;
  wire [2:0] _2950_;
  wire [2:0] _2951_;
  wire [2:0] _2952_;
  wire [2:0] _2953_;
  wire [2:0] _2954_;
  wire [2:0] _2955_;
  wire [2:0] _2956_;
  wire [2:0] _2957_;
  wire [2:0] _2958_;
  wire [2:0] _2959_;
  wire _2960_;
  wire [2:0] _2961_;
  wire [2:0] _2962_;
  wire [2:0] _2963_;
  wire _2964_;
  wire _2965_;
  wire [2:0] _2966_;
  wire [2:0] _2967_;
  wire [2:0] _2968_;
  wire [2:0] _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire [3:0] _2974_;
  wire [3:0] _2975_;
  wire [7:0] _2976_;
  wire [10:0] _2977_;
  wire [12:0] _2978_;
  wire [12:0] _2979_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3586" *)
  wire _2980_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _2981_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _2982_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _2983_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _2984_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _2985_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _2986_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _2987_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _2988_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3588" *)
  wire _2989_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _2990_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _2991_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _2992_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _2993_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _2994_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _2995_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _2996_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _2997_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3590" *)
  wire _2998_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _2999_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3000_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3001_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3002_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3003_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3004_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3005_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3006_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3592" *)
  wire _3007_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3008_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3009_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3010_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3011_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3012_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3013_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3014_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3015_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7781" *)
  wire _3016_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7784" *)
  wire _3017_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7785" *)
  wire _3018_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7786" *)
  wire _3019_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7787" *)
  wire _3020_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7788" *)
  wire _3021_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7789" *)
  wire _3022_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7790" *)
  wire _3023_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7791" *)
  wire _3024_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7952" *)
  wire _3025_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7953" *)
  wire _3026_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7954" *)
  wire _3027_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7955" *)
  wire _3028_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7956" *)
  wire _3029_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7957" *)
  wire _3030_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7958" *)
  wire _3031_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7959" *)
  wire _3032_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7960" *)
  wire _3033_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8787" *)
  wire _3034_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8850" *)
  wire _3035_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8851" *)
  wire _3036_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8852" *)
  wire _3037_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8853" *)
  wire _3038_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8854" *)
  wire _3039_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8855" *)
  wire _3040_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8856" *)
  wire _3041_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8857" *)
  wire _3042_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8910" *)
  wire _3043_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8911" *)
  wire _3044_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8912" *)
  wire _3045_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8913" *)
  wire _3046_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8922" *)
  wire _3047_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8923" *)
  wire _3048_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8924" *)
  wire _3049_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8925" *)
  wire _3050_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8926" *)
  wire _3051_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8927" *)
  wire _3052_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8928" *)
  wire _3053_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8929" *)
  wire _3054_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8983" *)
  wire _3055_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8984" *)
  wire _3056_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8985" *)
  wire _3057_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8986" *)
  wire _3058_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8994" *)
  wire _3059_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8995" *)
  wire _3060_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8996" *)
  wire _3061_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8997" *)
  wire _3062_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8998" *)
  wire _3063_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8999" *)
  wire _3064_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9000" *)
  wire _3065_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9001" *)
  wire _3066_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9099" *)
  wire _3067_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9100" *)
  wire _3068_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9101" *)
  wire _3069_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9102" *)
  wire _3070_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1186" *)
  wire _3071_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1189" *)
  wire [9:0] _3072_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1440" *)
  wire _3073_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3586" *)
  wire _3074_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _3075_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _3076_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _3077_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _3078_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _3079_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _3080_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _3081_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *)
  wire _3082_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3588" *)
  wire _3083_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _3084_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _3085_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _3086_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _3087_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _3088_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _3089_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _3090_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *)
  wire _3091_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3590" *)
  wire _3092_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3093_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3094_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3095_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3096_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3097_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3098_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3099_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *)
  wire _3100_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3592" *)
  wire _3101_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3102_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3103_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3104_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3105_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3106_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3107_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3108_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *)
  wire _3109_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4148" *)
  wire _3110_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5090" *)
  wire _3111_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5456" *)
  wire _3112_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5845" *)
  wire _3113_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6374" *)
  wire _3114_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6375" *)
  wire _3115_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6376" *)
  wire _3116_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6377" *)
  wire _3117_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6587" *)
  wire _3118_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6588" *)
  wire _3119_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6589" *)
  wire _3120_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6590" *)
  wire _3121_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6591" *)
  wire _3122_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6592" *)
  wire _3123_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6593" *)
  wire _3124_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6594" *)
  wire _3125_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7029" *)
  wire _3126_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7030" *)
  wire _3127_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7031" *)
  wire _3128_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7032" *)
  wire _3129_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7242" *)
  wire _3130_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7243" *)
  wire _3131_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7244" *)
  wire _3132_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7245" *)
  wire _3133_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7246" *)
  wire _3134_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7247" *)
  wire _3135_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7248" *)
  wire _3136_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7249" *)
  wire _3137_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8762" *)
  wire _3138_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1201" *)
  wire [31:0] _3139_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1451" *)
  wire [5:0] _3140_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1522" *)
  wire [2:0] _3141_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2175" *)
  wire [2:0] _3142_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3426" *)
  wire [31:0] _3143_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5841" *)
  wire [31:0] _3144_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1222" *)
  wire [12:0] _3145_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1222" *)
  wire [12:0] _3146_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2258" *)
  wire _3147_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3274" *)
  wire _3148_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3281" *)
  wire _3149_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3288" *)
  wire _3150_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3295" *)
  wire _3151_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3302" *)
  wire _3152_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3309" *)
  wire _3153_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3316" *)
  wire _3154_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3323" *)
  wire _3155_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3156_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3157_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3158_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3159_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3160_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3161_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3162_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3163_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3164_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3165_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3166_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3167_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3168_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3169_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3170_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3171_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3172_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3173_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3174_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3175_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3176_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3177_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3178_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3179_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3180_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3181_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3182_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3183_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3184_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3185_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3186_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *)
  wire [27:0] _3187_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3188_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3189_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3190_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3191_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3192_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3193_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3194_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3195_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3196_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3197_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3198_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3199_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3200_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3201_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3202_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3203_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3204_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3205_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3206_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3207_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3208_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3209_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3210_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3211_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3212_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3213_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3214_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3215_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3216_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3217_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3218_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *)
  wire [27:0] _3219_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3220_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3221_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3222_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3223_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3224_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3225_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3226_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3227_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3228_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3229_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3230_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3231_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3232_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3233_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3234_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3235_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3236_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3237_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3238_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3239_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3240_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3241_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3242_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3243_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3244_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3245_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3246_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3247_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3248_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3249_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3250_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3251_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3252_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3253_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3254_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3255_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3256_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3257_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3258_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3259_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3260_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3261_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3262_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3263_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3264_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3265_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3266_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3267_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3268_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3269_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3270_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3271_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3272_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3273_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3274_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3275_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3276_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3277_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3278_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3279_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3280_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3281_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3282_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *)
  wire [27:0] _3283_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3284_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3285_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3286_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3287_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3288_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3289_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3290_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3291_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3292_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3293_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3294_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3295_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3296_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3297_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3298_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3299_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3300_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3301_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3302_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3303_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3304_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3305_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3306_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3307_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3308_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3309_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3310_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3311_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3312_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3313_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3314_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *)
  wire [27:0] _3315_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3316_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3317_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3318_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3319_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3320_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3321_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3322_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3323_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3324_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3325_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3326_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3327_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3328_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3329_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3330_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3331_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3332_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3333_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3334_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3335_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3336_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3337_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3338_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3339_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3340_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3341_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3342_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3343_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3344_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3345_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3346_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3347_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3348_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3349_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3350_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3351_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3352_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3353_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3354_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3355_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3356_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3357_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3358_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3359_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3360_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3361_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3362_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3363_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3364_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3365_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3366_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3367_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3368_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3369_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3370_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3371_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3372_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3373_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3374_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3375_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3376_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3377_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3378_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *)
  wire [27:0] _3379_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3380_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3381_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3382_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3383_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3384_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3385_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3386_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3387_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3388_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3389_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3390_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3391_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3392_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3393_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3394_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3395_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3396_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3397_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3398_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3399_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3400_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3401_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3402_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3403_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3404_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3405_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3406_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3407_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3408_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3409_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3410_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *)
  wire [27:0] _3411_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [27:0] _3412_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [27:0] _3413_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [27:0] _3414_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [27:0] _3415_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [27:0] _3416_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [27:0] _3417_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [27:0] _3418_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *)
  wire [27:0] _3419_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3420_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3421_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3422_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3423_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3424_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3425_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3426_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3427_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3428_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3429_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3430_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3431_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3432_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3433_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3434_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *)
  wire [31:0] _3435_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [27:0] _3436_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [27:0] _3437_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [27:0] _3438_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [27:0] _3439_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [27:0] _3440_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [27:0] _3441_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [27:0] _3442_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *)
  wire [27:0] _3443_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3444_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3445_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3446_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3447_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3448_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3449_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3450_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3451_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3452_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3453_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3454_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3455_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3456_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3457_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *)
  wire [31:0] _3458_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [27:0] _3459_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [27:0] _3460_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [27:0] _3461_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [27:0] _3462_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [27:0] _3463_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [27:0] _3464_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [27:0] _3465_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *)
  wire [27:0] _3466_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3467_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3468_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3469_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3470_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3471_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3472_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3473_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3474_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3475_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3476_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3477_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3478_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3479_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3480_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3481_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *)
  wire [31:0] _3482_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [27:0] _3483_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [27:0] _3484_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [27:0] _3485_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [27:0] _3486_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [27:0] _3487_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [27:0] _3488_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [27:0] _3489_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *)
  wire [27:0] _3490_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _3491_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *)
  wire [31:0] _3492_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3645" *)
  wire [114:0] _3493_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3646" *)
  wire [114:0] _3494_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3647" *)
  wire [114:0] _3495_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3648" *)
  wire [114:0] _3496_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3649" *)
  wire [114:0] _3497_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3650" *)
  wire [114:0] _3498_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3651" *)
  wire [114:0] _3499_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3652" *)
  wire [114:0] _3500_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6386" *)
  wire [18:0] _3501_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6387" *)
  wire [18:0] _3502_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6388" *)
  wire [18:0] _3503_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6389" *)
  wire [18:0] _3504_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6611" *)
  wire [10:0] _3505_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6612" *)
  wire [10:0] _3506_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6613" *)
  wire [10:0] _3507_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6614" *)
  wire [10:0] _3508_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6615" *)
  wire [10:0] _3509_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6616" *)
  wire [10:0] _3510_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6617" *)
  wire [10:0] _3511_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6618" *)
  wire [10:0] _3512_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7041" *)
  wire [15:0] _3513_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7042" *)
  wire [15:0] _3514_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7043" *)
  wire [15:0] _3515_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7044" *)
  wire [15:0] _3516_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7266" *)
  wire [7:0] _3517_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7267" *)
  wire [7:0] _3518_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7268" *)
  wire [7:0] _3519_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7269" *)
  wire [7:0] _3520_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7270" *)
  wire [7:0] _3521_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7271" *)
  wire [7:0] _3522_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7272" *)
  wire [7:0] _3523_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7273" *)
  wire [7:0] _3524_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8023" *)
  wire [114:0] _3525_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8024" *)
  wire [114:0] _3526_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8025" *)
  wire [114:0] _3527_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8026" *)
  wire [114:0] _3528_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8027" *)
  wire [114:0] _3529_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8028" *)
  wire [114:0] _3530_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8029" *)
  wire [114:0] _3531_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8030" *)
  wire [114:0] _3532_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8031" *)
  wire [114:0] _3533_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8032" *)
  wire [114:0] _3534_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8033" *)
  wire [114:0] _3535_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8034" *)
  wire [114:0] _3536_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8035" *)
  wire [114:0] _3537_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8036" *)
  wire [114:0] _3538_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8037" *)
  wire [114:0] _3539_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8038" *)
  wire [114:0] _3540_;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:95" *)
  wire [5:0] BANK_DEPTH;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:96" *)
  wire active_last_line;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:97" *)
  wire average_pooling_en;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:746" *)
  wire [3:0] bank_merge_num;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:747" *)
  reg [2:0] bubble_add;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:748" *)
  reg [2:0] bubble_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:98" *)
  wire bubble_en_end;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:749" *)
  reg [2:0] bubble_num;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:99" *)
  wire [2:0] bubble_num_dec;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:750" *)
  reg [2:0] bubble_num_use;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:100" *)
  wire [3:0] buffer_lines_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:101" *)
  wire [3:0] buffer_lines_1;
  wire buffer_lines_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:103" *)
  wire [3:0] buffer_lines_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:751" *)
  reg [3:0] buffer_lines_num;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:752" *)
  reg [1:0] c_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:753" *)
  reg [1:0] channel_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:754" *)
  reg cube_end_flag;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:104" *)
  wire [3:0] cube_in_height_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:105" *)
  wire [13:0] cube_out_channel;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:755" *)
  reg cur_datin_disable;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:756" *)
  reg cur_datin_disable_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:106" *)
  wire cur_datin_disable_2d_sync;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:757" *)
  reg cur_datin_disable_3d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:758" *)
  reg cur_datin_disable_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:107" *)
  wire [21:0] data_16bit_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:108" *)
  wire [21:0] data_16bit_0_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:109" *)
  wire [21:0] data_16bit_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:110" *)
  wire [21:0] data_16bit_1_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:111" *)
  wire [21:0] data_16bit_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:112" *)
  wire [21:0] data_16bit_2_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:113" *)
  wire [21:0] data_16bit_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:114" *)
  wire [21:0] data_16bit_3_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:115" *)
  wire [13:0] data_8bit_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:116" *)
  wire [13:0] data_8bit_0_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:117" *)
  wire [13:0] data_8bit_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:118" *)
  wire [13:0] data_8bit_1_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:119" *)
  wire [13:0] data_8bit_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:120" *)
  wire [13:0] data_8bit_2_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:121" *)
  wire [13:0] data_8bit_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:122" *)
  wire [13:0] data_8bit_3_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:123" *)
  wire [13:0] data_8bit_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:124" *)
  wire [13:0] data_8bit_4_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:125" *)
  wire [13:0] data_8bit_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:126" *)
  wire [13:0] data_8bit_5_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:127" *)
  wire [13:0] data_8bit_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:128" *)
  wire [13:0] data_8bit_6_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:129" *)
  wire [13:0] data_8bit_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:130" *)
  wire [13:0] data_8bit_7_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:131" *)
  wire data_c_end;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:132" *)
  wire [18:0] data_hmult_16bit_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:133" *)
  (* unused_bits = "35 36 37" *)
  wire [38:0] data_hmult_16bit_0_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:134" *)
  wire [38:0] data_hmult_16bit_0_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:135" *)
  wire [18:0] data_hmult_16bit_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:136" *)
  (* unused_bits = "35 36 37" *)
  wire [38:0] data_hmult_16bit_1_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:137" *)
  wire [38:0] data_hmult_16bit_1_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:138" *)
  wire [18:0] data_hmult_16bit_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:139" *)
  (* unused_bits = "35 36 37" *)
  wire [38:0] data_hmult_16bit_2_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:140" *)
  wire [38:0] data_hmult_16bit_2_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:141" *)
  wire [18:0] data_hmult_16bit_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:142" *)
  (* unused_bits = "35 36 37" *)
  wire [38:0] data_hmult_16bit_3_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:143" *)
  wire [38:0] data_hmult_16bit_3_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:144" *)
  wire [21:0] data_hmult_8bit_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:145" *)
  (* unused_bits = "27 28 29" *)
  wire [30:0] data_hmult_8bit_0_lsb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:146" *)
  wire [30:0] data_hmult_8bit_0_lsb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:147" *)
  (* unused_bits = "27 28 29" *)
  wire [30:0] data_hmult_8bit_0_msb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:148" *)
  wire [30:0] data_hmult_8bit_0_msb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:149" *)
  wire [21:0] data_hmult_8bit_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:150" *)
  (* unused_bits = "27 28 29" *)
  wire [30:0] data_hmult_8bit_1_lsb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:151" *)
  wire [30:0] data_hmult_8bit_1_lsb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:152" *)
  (* unused_bits = "27 28 29" *)
  wire [30:0] data_hmult_8bit_1_msb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:153" *)
  wire [30:0] data_hmult_8bit_1_msb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:154" *)
  wire [21:0] data_hmult_8bit_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:155" *)
  (* unused_bits = "27 28 29" *)
  wire [30:0] data_hmult_8bit_2_lsb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:156" *)
  wire [30:0] data_hmult_8bit_2_lsb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:157" *)
  (* unused_bits = "27 28 29" *)
  wire [30:0] data_hmult_8bit_2_msb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:158" *)
  wire [30:0] data_hmult_8bit_2_msb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:159" *)
  wire [21:0] data_hmult_8bit_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:160" *)
  (* unused_bits = "27 28 29" *)
  wire [30:0] data_hmult_8bit_3_lsb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:161" *)
  wire [30:0] data_hmult_8bit_3_lsb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:162" *)
  (* unused_bits = "27 28 29" *)
  wire [30:0] data_hmult_8bit_3_msb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:163" *)
  wire [30:0] data_hmult_8bit_3_msb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:164" *)
  wire [21:0] data_hmult_stage0_in0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:165" *)
  wire [21:0] data_hmult_stage0_in1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:166" *)
  wire [21:0] data_hmult_stage0_in2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:167" *)
  wire [21:0] data_hmult_stage0_in3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:168" *)
  wire [15:0] data_mult_stage1_in0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:169" *)
  wire [15:0] data_mult_stage1_in1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:170" *)
  wire [15:0] data_mult_stage1_in2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:171" *)
  wire [15:0] data_mult_stage1_in3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:172" *)
  wire [15:0] data_vmult_16bit_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:173" *)
  (* unused_bits = "32 33 34" *)
  wire [35:0] data_vmult_16bit_0_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:174" *)
  wire [35:0] data_vmult_16bit_0_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:175" *)
  wire [15:0] data_vmult_16bit_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:176" *)
  (* unused_bits = "32 33 34" *)
  wire [35:0] data_vmult_16bit_1_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:177" *)
  wire [35:0] data_vmult_16bit_1_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:178" *)
  wire [15:0] data_vmult_16bit_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:179" *)
  (* unused_bits = "32 33 34" *)
  wire [35:0] data_vmult_16bit_2_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:180" *)
  wire [35:0] data_vmult_16bit_2_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:181" *)
  wire [15:0] data_vmult_16bit_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:182" *)
  (* unused_bits = "32 33 34" *)
  wire [35:0] data_vmult_16bit_3_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:183" *)
  wire [35:0] data_vmult_16bit_3_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:184" *)
  wire [15:0] data_vmult_8bit_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:185" *)
  (* unused_bits = "24 25 26" *)
  wire [27:0] data_vmult_8bit_0_lsb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:186" *)
  wire [27:0] data_vmult_8bit_0_lsb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:187" *)
  (* unused_bits = "24 25 26" *)
  wire [27:0] data_vmult_8bit_0_msb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:188" *)
  wire [27:0] data_vmult_8bit_0_msb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:189" *)
  wire [15:0] data_vmult_8bit_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:190" *)
  (* unused_bits = "24 25 26" *)
  wire [27:0] data_vmult_8bit_1_lsb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:191" *)
  wire [27:0] data_vmult_8bit_1_lsb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:192" *)
  (* unused_bits = "24 25 26" *)
  wire [27:0] data_vmult_8bit_1_msb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:193" *)
  wire [27:0] data_vmult_8bit_1_msb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:194" *)
  wire [15:0] data_vmult_8bit_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:195" *)
  (* unused_bits = "24 25 26" *)
  wire [27:0] data_vmult_8bit_2_lsb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:196" *)
  wire [27:0] data_vmult_8bit_2_lsb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:197" *)
  (* unused_bits = "24 25 26" *)
  wire [27:0] data_vmult_8bit_2_msb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:198" *)
  wire [27:0] data_vmult_8bit_2_msb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:199" *)
  wire [15:0] data_vmult_8bit_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:200" *)
  (* unused_bits = "24 25 26" *)
  wire [27:0] data_vmult_8bit_3_lsb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:201" *)
  wire [27:0] data_vmult_8bit_3_lsb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:202" *)
  (* unused_bits = "24 25 26" *)
  wire [27:0] data_vmult_8bit_3_msb_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:203" *)
  wire [27:0] data_vmult_8bit_3_msb_ext_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:759" *)
  reg [111:0] datin_buf;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:760" *)
  reg [111:0] datin_buf_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:204" *)
  wire [254:0] din_pd;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:205" *)
  wire [254:0] din_pd_d0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:206" *)
  wire [254:0] din_pd_d1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:207" *)
  wire [254:0] din_pd_d2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:208" *)
  wire [254:0] din_pd_d3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:209" *)
  wire [254:0] din_pd_d4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:210" *)
  wire din_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:211" *)
  wire din_rdy_d0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:212" *)
  wire din_rdy_d1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:213" *)
  wire din_rdy_d2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:214" *)
  wire din_rdy_d3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:215" *)
  wire din_rdy_d4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:216" *)
  wire din_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:217" *)
  wire din_vld_d0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:218" *)
  wire din_vld_d1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:219" *)
  wire din_vld_d2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:220" *)
  wire din_vld_d3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:221" *)
  wire din_vld_d4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:222" *)
  wire [254:0] dout_pd;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:223" *)
  wire dout_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:224" *)
  wire dout_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:225" *)
  wire [3:0] first_out_num;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:226" *)
  wire [2:0] first_out_num_dec2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:227" *)
  wire first_splitw;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:228" *)
  wire [2:0] flush_in_next_surf;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:761" *)
  wire [2:0] flush_num;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:762" *)
  wire [2:0] flush_num_cal;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:229" *)
  wire [2:0] flush_num_dec1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:230" *)
  wire flush_read_en;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:763" *)
  reg flush_read_en_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:231" *)
  wire [7:0] fp16_4add_in_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:232" *)
  wire [7:0] fp16_4add_in_pvld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:233" *)
  wire [7:0] fp16_4add_out_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:234" *)
  wire [7:0] fp16_4add_out_pvld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:235" *)
  wire [67:0] fp16_add_in_a;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:236" *)
  wire [67:0] fp16_add_in_a_sync;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:237" *)
  wire [67:0] fp16_add_in_b0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:238" *)
  wire [67:0] fp16_add_in_b1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:239" *)
  wire [67:0] fp16_add_in_b2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:240" *)
  wire [67:0] fp16_add_in_b3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:241" *)
  wire [67:0] fp16_add_in_b4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:242" *)
  wire [67:0] fp16_add_in_b5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:243" *)
  wire [67:0] fp16_add_in_b6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:244" *)
  wire [67:0] fp16_add_in_b7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:245" *)
  wire fp16_add_in_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:246" *)
  wire [3:0] fp16_add_pad_in_a_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:247" *)
  wire [3:0] fp16_add_pad_in_a_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:248" *)
  wire [3:0] fp16_add_pad_in_b_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:249" *)
  wire [3:0] fp16_add_pad_in_b_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:250" *)
  wire [16:0] fp16_add_pad_out0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:251" *)
  wire [16:0] fp16_add_pad_out1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:252" *)
  wire [16:0] fp16_add_pad_out2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:253" *)
  wire [16:0] fp16_add_pad_out3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:254" *)
  wire fp16_add_pad_out_pvld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:255" *)
  wire [3:0] fp16_add_pad_out_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:256" *)
  wire [3:0] fp16_add_pad_out_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:257" *)
  wire fp16_en;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:258" *)
  wire fp16_mean_pool_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:259" *)
  wire fp16_mean_pool_valid;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:260" *)
  wire [114:0] fp16_mul_pad_line_in_pd;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:261" *)
  wire [114:0] fp16_mul_pad_line_in_pd_d0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:262" *)
  wire [114:0] fp16_mul_pad_line_in_pd_d1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:263" *)
  wire [114:0] fp16_mul_pad_line_in_pd_d2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:264" *)
  wire [114:0] fp16_mul_pad_line_in_pd_d3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:265" *)
  wire fp16_mul_pad_line_in_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:266" *)
  wire fp16_mul_pad_line_in_rdy_d0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:267" *)
  wire fp16_mul_pad_line_in_rdy_d1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:268" *)
  wire fp16_mul_pad_line_in_rdy_d2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:269" *)
  wire fp16_mul_pad_line_in_rdy_d3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:270" *)
  wire fp16_mul_pad_line_in_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:271" *)
  wire fp16_mul_pad_line_in_vld_d0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:272" *)
  wire fp16_mul_pad_line_in_vld_d1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:273" *)
  wire fp16_mul_pad_line_in_vld_d2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:274" *)
  wire fp16_mul_pad_line_in_vld_d3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:275" *)
  wire [114:0] fp16_mul_pad_line_out_pd;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:276" *)
  wire fp16_mul_pad_line_out_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:277" *)
  wire fp16_mul_pad_line_out_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:278" *)
  wire fp16_mul_pad_line_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:279" *)
  wire fp16_mul_pad_line_pvld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:280" *)
  wire [1:0] fp16_mul_pad_line_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:281" *)
  wire [1:0] fp16_mul_pad_line_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:282" *)
  wire [3:0] fp16_mulv_in_a_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:283" *)
  wire [3:0] fp16_mulv_in_a_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:284" *)
  wire [3:0] fp16_mulv_in_b_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:285" *)
  wire [3:0] fp16_mulv_in_b_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:286" *)
  wire fp16_mulv_in_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:287" *)
  wire [16:0] fp16_mulv_out0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:288" *)
  wire [16:0] fp16_mulv_out1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:289" *)
  wire [16:0] fp16_mulv_out2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:290" *)
  wire [16:0] fp16_mulv_out3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:291" *)
  wire [3:0] fp16_mulv_out_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:292" *)
  wire [3:0] fp16_mulv_out_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:293" *)
  wire fp16_mulv_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:294" *)
  wire [3:0] fp16_mulw_in_a_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:295" *)
  wire [3:0] fp16_mulw_in_a_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:296" *)
  wire [3:0] fp16_mulw_in_b_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:297" *)
  wire [3:0] fp16_mulw_in_b_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:298" *)
  wire fp16_mulw_in_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:299" *)
  wire [16:0] fp16_mulw_out0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:300" *)
  wire [16:0] fp16_mulw_out1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:301" *)
  wire [16:0] fp16_mulw_out2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:302" *)
  wire [16:0] fp16_mulw_out3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:303" *)
  wire fp16_mulw_out_pvld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:304" *)
  wire [3:0] fp16_mulw_out_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:305" *)
  wire [3:0] fp16_mulw_out_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:306" *)
  wire fp16_mulw_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:307" *)
  wire [114:0] fp16_pout_mem_data;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:308" *)
  wire [15:0] fp17T16_out0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:309" *)
  wire [15:0] fp17T16_out1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:310" *)
  wire [15:0] fp17T16_out2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:311" *)
  wire [15:0] fp17T16_out3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:312" *)
  wire [3:0] fp17T16_out_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:313" *)
  wire [3:0] fp17T16_out_vld;
  wire [100:0] fp_add_out_dp_ext_0;
  wire [100:0] fp_add_out_dp_ext_1;
  wire [100:0] fp_add_out_dp_ext_2;
  wire [100:0] fp_add_out_dp_ext_3;
  wire [100:0] fp_add_out_dp_ext_4;
  wire [100:0] fp_add_out_dp_ext_5;
  wire [100:0] fp_add_out_dp_ext_6;
  wire [100:0] fp_add_out_dp_ext_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:322" *)
  wire fp_add_out_load;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:323" *)
  wire fp_add_out_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:324" *)
  wire [63:0] fp_dp2wdma_dp;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:325" *)
  wire fp_dp2wdma_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:326" *)
  wire fp_dp2wdma_pvld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:327" *)
  wire [5:0] fp_mem0_waddr;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:328" *)
  wire [115:0] fp_mem0_wdata;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:329" *)
  wire [5:0] fp_mem1_waddr;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:330" *)
  wire [115:0] fp_mem1_wdata;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:331" *)
  wire [5:0] fp_mem2_waddr;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:332" *)
  wire [115:0] fp_mem2_wdata;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:333" *)
  wire [5:0] fp_mem3_waddr;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:334" *)
  wire [115:0] fp_mem3_wdata;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:335" *)
  wire [5:0] fp_mem4_waddr;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:336" *)
  wire [115:0] fp_mem4_wdata;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:337" *)
  wire [5:0] fp_mem5_waddr;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:338" *)
  wire [115:0] fp_mem5_wdata;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:339" *)
  wire [5:0] fp_mem6_waddr;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:340" *)
  wire [115:0] fp_mem6_wdata;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:341" *)
  wire [5:0] fp_mem7_waddr;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:342" *)
  wire [115:0] fp_mem7_wdata;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:343" *)
  wire [2:0] fp_mem_size_v;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:344" *)
  wire [7:0] fp_mem_we;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:345" *)
  wire fp_mulw_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:346" *)
  wire [115:0] fp_pooling_result0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:347" *)
  wire [115:0] fp_pooling_result1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:348" *)
  wire [115:0] fp_pooling_result2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:349" *)
  wire [115:0] fp_pooling_result3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:350" *)
  wire [115:0] fp_pooling_result4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:351" *)
  wire [115:0] fp_pooling_result5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:352" *)
  wire [115:0] fp_pooling_result6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:353" *)
  wire [115:0] fp_pooling_result7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:354" *)
  wire [67:0] fp_pooling_result_dp_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:355" *)
  wire [67:0] fp_pooling_result_dp_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:356" *)
  wire [67:0] fp_pooling_result_dp_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:357" *)
  wire [67:0] fp_pooling_result_dp_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:358" *)
  wire [67:0] fp_pooling_result_dp_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:359" *)
  wire [67:0] fp_pooling_result_dp_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:360" *)
  wire [67:0] fp_pooling_result_dp_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:361" *)
  wire [67:0] fp_pooling_result_dp_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:362" *)
  wire [114:0] fp_pout_mem_data;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:363" *)
  wire [114:0] fp_pout_mem_data_act;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:364" *)
  wire [114:0] fp_pout_mem_data_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:365" *)
  wire [7:0] fp_pout_mem_data_sel;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:366" *)
  wire [7:0] fp_pout_mem_data_sel_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:367" *)
  wire [3:0] h_pt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:368" *)
  wire [4:0] h_pt_pb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:369" *)
  wire [10:0] hmult_8bit_0_lsb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:370" *)
  wire [10:0] hmult_8bit_0_msb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:371" *)
  wire [10:0] hmult_8bit_1_lsb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:372" *)
  wire [10:0] hmult_8bit_1_msb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:373" *)
  wire [10:0] hmult_8bit_2_lsb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:374" *)
  wire [10:0] hmult_8bit_2_msb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:375" *)
  wire [10:0] hmult_8bit_3_lsb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:376" *)
  wire [10:0] hmult_8bit_3_msb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:377" *)
  wire i16_less_neg_0_5_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:378" *)
  wire i16_less_neg_0_5_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:379" *)
  wire i16_less_neg_0_5_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:380" *)
  wire i16_less_neg_0_5_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:381" *)
  wire i16_more_neg_0_5_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:382" *)
  wire i16_more_neg_0_5_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:383" *)
  wire i16_more_neg_0_5_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:384" *)
  wire i16_more_neg_0_5_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:385" *)
  wire [18:0] i16_neg_add1_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:386" *)
  wire [18:0] i16_neg_add1_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:387" *)
  wire [18:0] i16_neg_add1_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:388" *)
  wire [18:0] i16_neg_add1_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:389" *)
  wire [15:0] i16_neg_vadd1_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:390" *)
  wire [15:0] i16_neg_vadd1_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:391" *)
  wire [15:0] i16_neg_vadd1_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:392" *)
  wire [15:0] i16_neg_vadd1_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:393" *)
  wire i16_vless_neg_0_5_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:394" *)
  wire i16_vless_neg_0_5_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:395" *)
  wire i16_vless_neg_0_5_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:396" *)
  wire i16_vless_neg_0_5_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:397" *)
  wire i16_vmore_neg_0_5_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:398" *)
  wire i16_vmore_neg_0_5_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:399" *)
  wire i16_vmore_neg_0_5_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:400" *)
  wire i16_vmore_neg_0_5_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:401" *)
  wire i8_less_neg_0_5_0_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:402" *)
  wire i8_less_neg_0_5_0_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:403" *)
  wire i8_less_neg_0_5_1_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:404" *)
  wire i8_less_neg_0_5_1_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:405" *)
  wire i8_less_neg_0_5_2_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:406" *)
  wire i8_less_neg_0_5_2_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:407" *)
  wire i8_less_neg_0_5_3_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:408" *)
  wire i8_less_neg_0_5_3_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:409" *)
  wire i8_more_neg_0_5_0_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:410" *)
  wire i8_more_neg_0_5_0_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:411" *)
  wire i8_more_neg_0_5_1_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:412" *)
  wire i8_more_neg_0_5_1_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:413" *)
  wire i8_more_neg_0_5_2_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:414" *)
  wire i8_more_neg_0_5_2_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:415" *)
  wire i8_more_neg_0_5_3_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:416" *)
  wire i8_more_neg_0_5_3_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:417" *)
  wire [10:0] i8_neg_add1_0_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:418" *)
  wire [10:0] i8_neg_add1_0_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:419" *)
  wire [10:0] i8_neg_add1_1_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:420" *)
  wire [10:0] i8_neg_add1_1_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:421" *)
  wire [10:0] i8_neg_add1_2_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:422" *)
  wire [10:0] i8_neg_add1_2_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:423" *)
  wire [10:0] i8_neg_add1_3_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:424" *)
  wire [10:0] i8_neg_add1_3_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:425" *)
  wire [7:0] i8_neg_vadd1_0_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:426" *)
  wire [7:0] i8_neg_vadd1_0_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:427" *)
  wire [7:0] i8_neg_vadd1_1_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:428" *)
  wire [7:0] i8_neg_vadd1_1_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:429" *)
  wire [7:0] i8_neg_vadd1_2_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:430" *)
  wire [7:0] i8_neg_vadd1_2_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:431" *)
  wire [7:0] i8_neg_vadd1_3_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:432" *)
  wire [7:0] i8_neg_vadd1_3_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:433" *)
  wire i8_vless_neg_0_5_0_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:434" *)
  wire i8_vless_neg_0_5_0_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:435" *)
  wire i8_vless_neg_0_5_1_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:436" *)
  wire i8_vless_neg_0_5_1_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:437" *)
  wire i8_vless_neg_0_5_2_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:438" *)
  wire i8_vless_neg_0_5_2_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:439" *)
  wire i8_vless_neg_0_5_3_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:440" *)
  wire i8_vless_neg_0_5_3_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:441" *)
  wire i8_vmore_neg_0_5_0_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:442" *)
  wire i8_vmore_neg_0_5_0_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:443" *)
  wire i8_vmore_neg_0_5_1_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:444" *)
  wire i8_vmore_neg_0_5_1_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:445" *)
  wire i8_vmore_neg_0_5_2_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:446" *)
  wire i8_vmore_neg_0_5_2_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:447" *)
  wire i8_vmore_neg_0_5_3_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:448" *)
  wire i8_vmore_neg_0_5_3_m;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:449" *)
  wire init_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:450" *)
  wire [7:0] init_unit2d_set;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:452" *)
  wire int8_en;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:453" *)
  wire [63:0] int_dp2wdma_pd;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:454" *)
  wire int_dp2wdma_valid;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:764" *)
  reg [5:0] int_mem_waddr;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:765" *)
  reg [115:0] int_mem_wdata_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:766" *)
  reg [115:0] int_mem_wdata_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:767" *)
  reg [115:0] int_mem_wdata_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:768" *)
  reg [115:0] int_mem_wdata_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:769" *)
  reg [115:0] int_mem_wdata_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:770" *)
  reg [115:0] int_mem_wdata_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:771" *)
  reg [115:0] int_mem_wdata_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:772" *)
  reg [115:0] int_mem_wdata_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:773" *)
  reg [7:0] int_mem_we;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:455" *)
  wire [114:0] int_pout_mem_data;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:774" *)
  wire is_one_width_in;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:456" *)
  wire [3:0] kernel_width_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:775" *)
  wire [16:0] kernel_width_fp17;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:776" *)
  reg last_active_line_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:777" *)
  reg last_active_line_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:457" *)
  wire last_c;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:458" *)
  wire last_line_in;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:778" *)
  reg [2:0] last_out_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:459" *)
  wire last_out_done;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:779" *)
  reg last_out_en;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:460" *)
  wire last_pooling_flag;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:461" *)
  wire last_splitw;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:462" *)
  wire last_sub_lbuf_done;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:780" *)
  reg [12:0] line_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:463" *)
  wire line_end;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:464" *)
  wire load_din;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:465" *)
  wire load_din_all;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:466" *)
  wire load_wr_stage1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:467" *)
  wire load_wr_stage1_all;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:468" *)
  wire load_wr_stage2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:469" *)
  wire load_wr_stage2_all;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:470" *)
  wire load_wr_stage3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:471" *)
  wire load_wr_stage3_all;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:781" *)
  reg [114:0] mem_data0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:782" *)
  reg [114:0] mem_data0_lst;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:783" *)
  reg [114:0] mem_data1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:784" *)
  reg [114:0] mem_data1_lst;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:785" *)
  reg [114:0] mem_data2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:786" *)
  reg [114:0] mem_data2_lst;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:787" *)
  reg [114:0] mem_data3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:788" *)
  reg [114:0] mem_data3_lst;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:789" *)
  reg [114:0] mem_data4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:790" *)
  reg [114:0] mem_data4_lst;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:791" *)
  reg [114:0] mem_data5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:792" *)
  reg [114:0] mem_data5_lst;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:793" *)
  reg [114:0] mem_data6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:794" *)
  reg [114:0] mem_data6_lst;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:795" *)
  reg [114:0] mem_data7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:796" *)
  reg [114:0] mem_data7_lst;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:472" *)
  wire [7:0] mem_data_valid;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:473" *)
  wire [5:0] mem_raddr;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:797" *)
  reg [5:0] mem_raddr_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:474" *)
  wire [5:0] mem_raddr_2d_sync;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:798" *)
  reg [5:0] mem_raddr_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:475" *)
  (* unused_bits = "115" *)
  wire [115:0] mem_rdata_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:476" *)
  (* unused_bits = "115" *)
  wire [115:0] mem_rdata_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:477" *)
  (* unused_bits = "115" *)
  wire [115:0] mem_rdata_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:478" *)
  (* unused_bits = "115" *)
  wire [115:0] mem_rdata_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:479" *)
  (* unused_bits = "115" *)
  wire [115:0] mem_rdata_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:480" *)
  (* unused_bits = "115" *)
  wire [115:0] mem_rdata_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:481" *)
  (* unused_bits = "115" *)
  wire [115:0] mem_rdata_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:482" *)
  (* unused_bits = "115" *)
  wire [115:0] mem_rdata_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:483" *)
  wire [7:0] mem_re;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:484" *)
  wire [7:0] mem_re1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:485" *)
  wire [7:0] mem_re1_1st;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:799" *)
  reg mem_re1_sel;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:486" *)
  wire [7:0] mem_re2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:487" *)
  wire [7:0] mem_re2_1st;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:488" *)
  wire [7:0] mem_re2_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:800" *)
  reg mem_re2_sel;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:801" *)
  reg mem_re2_sel_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:489" *)
  wire [7:0] mem_re3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:490" *)
  wire [7:0] mem_re3_1st;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:491" *)
  wire [7:0] mem_re3_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:802" *)
  reg mem_re3_sel;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:803" *)
  reg mem_re3_sel_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:492" *)
  wire [7:0] mem_re4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:493" *)
  wire [7:0] mem_re4_1st;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:494" *)
  wire [7:0] mem_re4_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:804" *)
  reg mem_re4_sel;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:805" *)
  reg mem_re4_sel_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:495" *)
  wire [7:0] mem_re_1st;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:806" *)
  reg [7:0] mem_re_1st_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:496" *)
  wire [7:0] mem_re_1st_2d_sync;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:807" *)
  reg [7:0] mem_re_1st_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:808" *)
  reg [7:0] mem_re_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:497" *)
  wire [7:0] mem_re_2d_sync;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:809" *)
  reg [7:0] mem_re_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:498" *)
  wire [7:0] mem_re_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:810" *)
  reg [7:0] mem_re_last_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:811" *)
  reg [7:0] mem_re_last_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:499" *)
  wire [5:0] mem_waddr_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:500" *)
  wire [5:0] mem_waddr_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:501" *)
  wire [5:0] mem_waddr_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:502" *)
  wire [5:0] mem_waddr_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:503" *)
  wire [5:0] mem_waddr_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:504" *)
  wire [5:0] mem_waddr_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:505" *)
  wire [5:0] mem_waddr_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:506" *)
  wire [5:0] mem_waddr_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:507" *)
  wire [115:0] mem_wdata_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:508" *)
  wire [115:0] mem_wdata_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:509" *)
  wire [115:0] mem_wdata_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:510" *)
  wire [115:0] mem_wdata_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:511" *)
  wire [115:0] mem_wdata_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:512" *)
  wire [115:0] mem_wdata_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:513" *)
  wire [115:0] mem_wdata_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:514" *)
  wire [115:0] mem_wdata_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:515" *)
  wire [7:0] mem_we;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:516" *)
  wire middle_surface_trig;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:517" *)
  wire mon_data_16bit_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:519" *)
  wire mon_data_16bit_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:521" *)
  wire mon_data_16bit_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:523" *)
  wire mon_data_16bit_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:525" *)
  wire [1:0] mon_data_8bit_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:526" *)
  (* unused_bits = "0 1" *)
  wire [1:0] mon_data_8bit_0_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:527" *)
  wire [1:0] mon_data_8bit_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:528" *)
  (* unused_bits = "0 1" *)
  wire [1:0] mon_data_8bit_1_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:529" *)
  wire [1:0] mon_data_8bit_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:530" *)
  (* unused_bits = "0 1" *)
  wire [1:0] mon_data_8bit_2_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:531" *)
  wire [1:0] mon_data_8bit_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:532" *)
  (* unused_bits = "0 1" *)
  wire [1:0] mon_data_8bit_3_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:533" *)
  wire [1:0] mon_data_8bit_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:534" *)
  (* unused_bits = "0 1" *)
  wire [1:0] mon_data_8bit_4_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:535" *)
  wire [1:0] mon_data_8bit_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:536" *)
  (* unused_bits = "0 1" *)
  wire [1:0] mon_data_8bit_5_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:537" *)
  wire [1:0] mon_data_8bit_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:538" *)
  (* unused_bits = "0 1" *)
  wire [1:0] mon_data_8bit_6_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:539" *)
  wire [1:0] mon_data_8bit_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:540" *)
  (* unused_bits = "0 1" *)
  wire [1:0] mon_data_8bit_7_ff;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:541" *)
  wire mon_first_out_num;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:812" *)
  reg need_bubble;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:575" *)
  wire need_flush;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:813" *)
  wire [2:0] next2_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:814" *)
  wire [2:0] next2_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:815" *)
  wire [2:0] next3_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:816" *)
  wire [2:0] next3_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:817" *)
  wire [2:0] next3_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:818" *)
  wire [2:0] next4_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:819" *)
  wire [2:0] next4_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:820" *)
  wire [2:0] next4_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:821" *)
  wire [2:0] next4_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:822" *)
  wire [2:0] next5_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:823" *)
  wire [2:0] next5_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:824" *)
  wire [2:0] next5_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:825" *)
  wire [2:0] next5_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:826" *)
  wire [2:0] next5_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:827" *)
  wire [2:0] next6_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:828" *)
  wire [2:0] next6_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:829" *)
  wire [2:0] next6_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:830" *)
  wire [2:0] next6_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:831" *)
  wire [2:0] next6_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:832" *)
  wire [2:0] next6_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:833" *)
  wire [2:0] next7_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:834" *)
  wire [2:0] next7_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:835" *)
  wire [2:0] next7_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:836" *)
  wire [2:0] next7_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:837" *)
  wire [2:0] next7_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:838" *)
  wire [2:0] next7_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:839" *)
  wire [2:0] next7_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:53" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:54" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:55" *)
  input nvdla_op_gated_clk_fp16;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:840" *)
  reg [2:0] one_width_bubble_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:576" *)
  wire one_width_bubble_end;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:841" *)
  reg one_width_disable;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:842" *)
  reg one_width_disable_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:577" *)
  wire one_width_disable_2d_sync;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:843" *)
  reg one_width_disable_3d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:844" *)
  reg one_width_disable_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:578" *)
  wire one_width_norm_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:579" *)
  wire [2:0] pad_l;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:580" *)
  wire [16:0] pad_line_sum;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:581" *)
  wire pad_line_sum_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:582" *)
  wire pad_line_sum_pvld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:583" *)
  wire [2:0] pad_r;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:845" *)
  wire [5:0] pad_r_remain;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:584" *)
  wire [2:0] pad_table_index;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:846" *)
  wire [18:0] pad_table_out;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:585" *)
  wire [21:0] pad_value;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:586" *)
  wire padding_here;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:587" *)
  wire [2:0] padding_stride1_num;
  wire [1:0] padding_stride2_num;
  wire [1:0] padding_stride3_num;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:590" *)
  wire [2:0] padding_stride4_num;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:847" *)
  wire [2:0] padding_stride_num;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:56" *)
  input [2:0] padding_v_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:92" *)
  output [63:0] pdp_dp2wdma_pd;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:57" *)
  input pdp_dp2wdma_ready;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:93" *)
  output pdp_dp2wdma_valid;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:58" *)
  input pdp_op_start;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:848" *)
  reg [2:0] pnum_flush0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:849" *)
  reg [2:0] pnum_flush1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:850" *)
  reg [2:0] pnum_flush2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:851" *)
  reg [2:0] pnum_flush3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:852" *)
  reg [2:0] pnum_flush4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:853" *)
  reg [2:0] pnum_flush5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:854" *)
  reg [2:0] pnum_flush6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:591" *)
  wire pooling1d_norm_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:59" *)
  input [111:0] pooling1d_pd;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:592" *)
  wire [111:0] pooling1d_pd_use;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:94" *)
  output pooling1d_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:593" *)
  wire pooling1d_prdy_use;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:60" *)
  input pooling1d_pvld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:594" *)
  wire pooling1d_pvld_use;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:595" *)
  wire pooling1d_vld_rebuild;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:596" *)
  wire [31:0] pooling_2d_info;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:597" *)
  wire [3:0] pooling_2d_info_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:598" *)
  wire [3:0] pooling_2d_info_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:599" *)
  wire [3:0] pooling_2d_info_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:600" *)
  wire [3:0] pooling_2d_info_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:601" *)
  wire [3:0] pooling_2d_info_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:602" *)
  wire [3:0] pooling_2d_info_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:603" *)
  wire [3:0] pooling_2d_info_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:604" *)
  wire [3:0] pooling_2d_info_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:605" *)
  wire [31:0] pooling_2d_info_sync;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:606" *)
  wire pooling_2d_rdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:607" *)
  wire [111:0] pooling_2d_result_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:608" *)
  wire [111:0] pooling_2d_result_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:609" *)
  wire [111:0] pooling_2d_result_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:610" *)
  wire [111:0] pooling_2d_result_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:611" *)
  wire [111:0] pooling_2d_result_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:612" *)
  wire [111:0] pooling_2d_result_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:613" *)
  wire [111:0] pooling_2d_result_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:614" *)
  wire [111:0] pooling_2d_result_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:61" *)
  input [12:0] pooling_channel_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:615" *)
  wire [111:0] pooling_datin;
  wire [100:0] pooling_datin_ext;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:62" *)
  input [9:0] pooling_out_fwidth_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:63" *)
  input [9:0] pooling_out_lwidth_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:64" *)
  input [9:0] pooling_out_mwidth_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:617" *)
  wire [3:0] pooling_size;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:618" *)
  wire [2:0] pooling_size_minus_sride;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:619" *)
  wire [3:0] pooling_size_v;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:65" *)
  input [2:0] pooling_size_v_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:66" *)
  input [7:0] pooling_splitw_num_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:620" *)
  wire pooling_stride_big;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:621" *)
  wire [4:0] pooling_stride_v;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:67" *)
  input [3:0] pooling_stride_v_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:68" *)
  input [1:0] pooling_type_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:855" *)
  reg [27:0] pout_data_0_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:856" *)
  reg [27:0] pout_data_0_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:857" *)
  reg [27:0] pout_data_0_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:858" *)
  reg [27:0] pout_data_0_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:859" *)
  reg [21:0] pout_data_stage0_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:860" *)
  reg [21:0] pout_data_stage0_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:861" *)
  reg [21:0] pout_data_stage0_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:862" *)
  reg [21:0] pout_data_stage0_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:622" *)
  wire pout_data_stage0_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:863" *)
  reg [15:0] pout_data_stage1_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:864" *)
  reg [15:0] pout_data_stage1_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:865" *)
  reg [15:0] pout_data_stage1_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:866" *)
  reg [15:0] pout_data_stage1_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:623" *)
  wire pout_data_stage1_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:867" *)
  reg pout_data_stage1_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:624" *)
  wire pout_data_stage2_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:868" *)
  reg pout_data_stage2_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:625" *)
  wire pout_data_stage3_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:869" *)
  reg pout_data_stage3_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:626" *)
  wire [114:0] pout_mem_data;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:627" *)
  wire [21:0] pout_mem_data0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:628" *)
  wire [21:0] pout_mem_data1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:629" *)
  wire [21:0] pout_mem_data2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:630" *)
  wire [21:0] pout_mem_data3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:870" *)
  reg [27:0] pout_mem_data_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:871" *)
  reg [27:0] pout_mem_data_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:872" *)
  reg [27:0] pout_mem_data_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:873" *)
  reg [27:0] pout_mem_data_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:874" *)
  wire [114:0] pout_mem_data_act;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:631" *)
  wire [114:0] pout_mem_data_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:632" *)
  wire [114:0] pout_mem_data_last_sync;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:633" *)
  wire [7:0] pout_mem_data_sel;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:634" *)
  wire [7:0] pout_mem_data_sel_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:635" *)
  wire [7:0] pout_mem_data_sel_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:636" *)
  wire [7:0] pout_mem_data_sel_1_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:637" *)
  wire [7:0] pout_mem_data_sel_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:638" *)
  wire [7:0] pout_mem_data_sel_2_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:639" *)
  wire [7:0] pout_mem_data_sel_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:640" *)
  wire [7:0] pout_mem_data_sel_3_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:641" *)
  wire [7:0] pout_mem_data_sel_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:642" *)
  wire [7:0] pout_mem_data_sel_last_sync;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:643" *)
  wire [7:0] pout_mem_data_sel_sync;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:875" *)
  reg [2:0] pout_mem_size_v;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:644" *)
  wire [2:0] pout_mem_size_v_use;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:645" *)
  wire [12:0] pout_width_cur;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:876" *)
  reg [12:0] pout_width_cur_latch;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:69" *)
  input [31:0] pwrbus_ram_pd;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:877" *)
  reg [2:0] rd_comb_lbuf_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:646" *)
  wire rd_comb_lbuf_end;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:647" *)
  wire rd_lbuf_end;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:648" *)
  wire rd_line_out;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:878" *)
  reg [5:0] rd_line_out_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:649" *)
  wire rd_line_out_done;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:650" *)
  wire rd_pout_data_en;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:879" *)
  reg rd_pout_data_en_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:880" *)
  reg rd_pout_data_en_3d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:881" *)
  reg rd_pout_data_en_4d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:882" *)
  reg rd_pout_data_en_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:651" *)
  wire rd_pout_data_stage0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:652" *)
  wire rd_pout_data_stage1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:653" *)
  wire rd_pout_data_stage1_all;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:654" *)
  wire rd_pout_data_stage2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:655" *)
  wire rd_pout_data_stage2_all;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:883" *)
  reg [2:0] rd_sub_lbuf_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:656" *)
  wire rd_sub_lbuf_end;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:70" *)
  input [12:0] reg2dp_cube_in_height;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:71" *)
  input [12:0] reg2dp_cube_out_width;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:72" *)
  input reg2dp_fp16_en;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:73" *)
  input [1:0] reg2dp_input_data;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:74" *)
  input reg2dp_int16_en;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:75" *)
  input reg2dp_int8_en;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:76" *)
  input [2:0] reg2dp_kernel_height;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:77" *)
  input [2:0] reg2dp_kernel_width;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:78" *)
  input [2:0] reg2dp_pad_bottom_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:79" *)
  input [2:0] reg2dp_pad_top;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:80" *)
  input [18:0] reg2dp_pad_value_1x_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:81" *)
  input [18:0] reg2dp_pad_value_2x_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:82" *)
  input [18:0] reg2dp_pad_value_3x_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:83" *)
  input [18:0] reg2dp_pad_value_4x_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:84" *)
  input [18:0] reg2dp_pad_value_5x_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:85" *)
  input [18:0] reg2dp_pad_value_6x_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:86" *)
  input [18:0] reg2dp_pad_value_7x_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:87" *)
  input [9:0] reg2dp_partial_width_out_first;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:88" *)
  input [9:0] reg2dp_partial_width_out_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:89" *)
  input [9:0] reg2dp_partial_width_out_mid;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:90" *)
  input [16:0] reg2dp_recip_height_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:884" *)
  reg [16:0] reg2dp_recip_height_use;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:91" *)
  input [16:0] reg2dp_recip_width_cfg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:885" *)
  reg [16:0] reg2dp_recip_width_use;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:657" *)
  wire [12:0] rest_height;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:658" *)
  wire [13:0] rest_height_use;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:886" *)
  wire [2:0] samllH_flush_num;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:659" *)
  wire small_active;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:660" *)
  wire splitw_enable;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:661" *)
  wire [4:0] stride;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:662" *)
  wire [4:0] stride_1x;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:663" *)
  wire [5:0] stride_2x;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:664" *)
  wire [6:0] stride_3x;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:665" *)
  wire [6:0] stride_4x;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:666" *)
  wire [7:0] stride_5x;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:667" *)
  wire [7:0] stride_6x;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:668" *)
  wire [7:0] stride_7x;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:669" *)
  wire stride_end;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:670" *)
  wire stride_trig_end;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:671" *)
  wire [2:0] strip_ycnt_offset;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:887" *)
  reg [2:0] strip_ycnt_psize;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:888" *)
  reg [3:0] strip_ycnt_stride;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:889" *)
  wire [3:0] strip_ycnt_stride_f;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:672" *)
  wire stripe_receive_done;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:890" *)
  reg [5:0] sub_lbuf_dout_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:673" *)
  wire sub_lbuf_dout_done;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:891" *)
  reg subend_need_flush_flg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:892" *)
  reg [10:0] surface_cnt_rd;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:674" *)
  wire [9:0] surface_num;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:675" *)
  wire [9:0] surface_num_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:676" *)
  wire [9:0] surface_num_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:893" *)
  reg surfend_need_bubble_flg;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:677" *)
  wire [7:0] unit2d_clr;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:894" *)
  reg [2:0] unit2d_cnt_pooling;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:678" *)
  wire [3:0] unit2d_cnt_pooling_a1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:679" *)
  wire [3:0] unit2d_cnt_pooling_a2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:680" *)
  wire [3:0] unit2d_cnt_pooling_a3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:681" *)
  wire [3:0] unit2d_cnt_pooling_a4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:682" *)
  wire [3:0] unit2d_cnt_pooling_a5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:683" *)
  wire [3:0] unit2d_cnt_pooling_a6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:684" *)
  wire [3:0] unit2d_cnt_pooling_a7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:685" *)
  wire unit2d_cnt_pooling_end;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:895" *)
  reg [2:0] unit2d_cnt_pooling_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:896" *)
  reg [2:0] unit2d_cnt_pooling_last_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:897" *)
  reg [2:0] unit2d_cnt_pooling_last_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:686" *)
  wire unit2d_cnt_pooling_last_end;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:687" *)
  wire [2:0] unit2d_cnt_pooling_max;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:898" *)
  reg [2:0] unit2d_cnt_stride;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:899" *)
  reg [7:0] unit2d_en;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:688" *)
  wire [7:0] unit2d_en_last;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:900" *)
  reg [7:0] unit2d_mem_1strd;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:689" *)
  wire [7:0] unit2d_set;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:690" *)
  wire [7:0] unit2d_set_trig;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:691" *)
  wire [2:0] unit2d_vsize1_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:692" *)
  wire [2:0] unit2d_vsize1_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:693" *)
  wire [2:0] unit2d_vsize1_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:694" *)
  wire [2:0] unit2d_vsize1_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:695" *)
  wire [2:0] unit2d_vsize1_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:696" *)
  wire [2:0] unit2d_vsize1_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:697" *)
  wire [2:0] unit2d_vsize1_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:698" *)
  wire [2:0] unit2d_vsize1_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:699" *)
  wire [2:0] unit2d_vsize2_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:700" *)
  wire [2:0] unit2d_vsize2_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:701" *)
  wire [2:0] unit2d_vsize2_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:702" *)
  wire [2:0] unit2d_vsize2_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:703" *)
  wire [2:0] unit2d_vsize2_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:704" *)
  wire [2:0] unit2d_vsize2_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:705" *)
  wire [2:0] unit2d_vsize2_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:706" *)
  wire [2:0] unit2d_vsize2_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:707" *)
  wire [2:0] unit2d_vsize3_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:708" *)
  wire [2:0] unit2d_vsize3_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:709" *)
  wire [2:0] unit2d_vsize3_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:710" *)
  wire [2:0] unit2d_vsize3_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:711" *)
  wire [2:0] unit2d_vsize3_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:712" *)
  wire [2:0] unit2d_vsize3_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:713" *)
  wire [2:0] unit2d_vsize3_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:714" *)
  wire [2:0] unit2d_vsize3_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:715" *)
  wire [2:0] unit2d_vsize4_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:716" *)
  wire [2:0] unit2d_vsize4_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:717" *)
  wire [2:0] unit2d_vsize4_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:718" *)
  wire [2:0] unit2d_vsize4_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:719" *)
  wire [2:0] unit2d_vsize4_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:720" *)
  wire [2:0] unit2d_vsize4_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:721" *)
  wire [2:0] unit2d_vsize4_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:722" *)
  wire [2:0] unit2d_vsize4_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:723" *)
  wire [2:0] unit2d_vsize_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:724" *)
  wire [2:0] unit2d_vsize_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:725" *)
  wire [2:0] unit2d_vsize_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:726" *)
  wire [2:0] unit2d_vsize_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:727" *)
  wire [2:0] unit2d_vsize_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:728" *)
  wire [2:0] unit2d_vsize_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:729" *)
  wire [2:0] unit2d_vsize_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:730" *)
  wire [2:0] unit2d_vsize_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:901" *)
  reg [2:0] unit2d_vsize_cnt_0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:902" *)
  reg [2:0] unit2d_vsize_cnt_0_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:903" *)
  reg [2:0] unit2d_vsize_cnt_1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:904" *)
  reg [2:0] unit2d_vsize_cnt_1_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:905" *)
  reg [2:0] unit2d_vsize_cnt_2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:906" *)
  reg [2:0] unit2d_vsize_cnt_2_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:907" *)
  reg [2:0] unit2d_vsize_cnt_3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:908" *)
  reg [2:0] unit2d_vsize_cnt_3_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:909" *)
  reg [2:0] unit2d_vsize_cnt_4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:910" *)
  reg [2:0] unit2d_vsize_cnt_4_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:911" *)
  reg [2:0] unit2d_vsize_cnt_5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:912" *)
  reg [2:0] unit2d_vsize_cnt_5_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:913" *)
  reg [2:0] unit2d_vsize_cnt_6;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:914" *)
  reg [2:0] unit2d_vsize_cnt_6_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:915" *)
  reg [2:0] unit2d_vsize_cnt_7;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:916" *)
  reg [2:0] unit2d_vsize_cnt_7_d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:731" *)
  wire [2:0] up_pnum0;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:917" *)
  reg up_pnum1;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:918" *)
  reg [1:0] up_pnum2;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:919" *)
  reg [1:0] up_pnum3;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:920" *)
  reg [2:0] up_pnum4;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:921" *)
  reg [2:0] up_pnum5;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:732" *)
  wire [7:0] vmult_8bit_0_lsb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:733" *)
  wire [7:0] vmult_8bit_0_msb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:734" *)
  wire [7:0] vmult_8bit_1_lsb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:735" *)
  wire [7:0] vmult_8bit_1_msb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:736" *)
  wire [7:0] vmult_8bit_2_lsb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:737" *)
  wire [7:0] vmult_8bit_2_msb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:738" *)
  wire [7:0] vmult_8bit_3_lsb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:739" *)
  wire [7:0] vmult_8bit_3_msb;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:740" *)
  wire wr_data_stage0_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:922" *)
  reg wr_data_stage0_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:741" *)
  wire wr_data_stage1_prdy;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:923" *)
  reg wr_data_stage1_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:924" *)
  reg wr_data_stage2_vld;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:925" *)
  reg [12:0] wr_line_dat_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:742" *)
  wire wr_line_dat_done;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:926" *)
  reg wr_line_end_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:927" *)
  reg wr_line_end_buf;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:928" *)
  reg [7:0] wr_splitc_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:929" *)
  reg [2:0] wr_sub_lbuf_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:743" *)
  wire wr_subcube_dat_done;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:930" *)
  reg [12:0] wr_surface_dat_cnt;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:744" *)
  wire wr_surface_dat_done;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:931" *)
  reg wr_surface_dat_done_2d;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:932" *)
  reg wr_surface_dat_done_buf;
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:745" *)
  wire wr_total_cube_done;
  assign _1230_ = c_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1153" *) 1'b1;
  assign _1231_ = wr_line_dat_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1165" *) 1'b1;
  assign _1232_ = wr_surface_dat_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1177" *) 1'b1;
  assign cube_out_channel = pooling_channel_cfg + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1183" *) 1'b1;
  assign surface_num_0 = cube_out_channel[13:4] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1186" *) _3071_;
  assign surface_num_1 = cube_out_channel[13:5] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1189" *) _3072_[0];
  assign _1233_[10:0] = surface_cnt_rd + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1198" *) 1'b1;
  assign _1234_ = wr_splitc_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1210" *) 1'b1;
  assign buffer_lines_1 = buffer_lines_0[3:1] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1234" *) buffer_lines_0[0];
  assign pooling_stride_v = pooling_stride_v_cfg + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1283" *) 1'b1;
  assign _1235_ = strip_ycnt_stride + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1317" *) 1'b1;
  assign _1236_[2:0] = strip_ycnt_psize + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1394" *) 1'b1;
  assign buffer_lines_0 = pooling_size_v_cfg + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1404" *) 1'b1;
  assign h_pt = reg2dp_cube_in_height[2:0] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1440" *) reg2dp_pad_top;
  assign h_pt_pb = h_pt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1443" *) reg2dp_pad_bottom_cfg;
  assign stride_3x = { pooling_stride_v, 1'b0 } + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1496" *) pooling_stride_v;
  assign stride_5x = { pooling_stride_v, 2'b00 } + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1498" *) pooling_stride_v;
  assign stride_6x = stride_3x + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1499" *) stride_3x;
  assign stride_7x = { pooling_stride_v, 2'b00 } + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1500" *) stride_3x;
  assign cube_in_height_cfg = reg2dp_cube_in_height[2:0] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1503" *) 1'b1;
  assign _1237_ = _3141_ + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1522" *) 1'b1;
  assign _1238_ = _1237_ + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1522" *) bubble_add;
  assign unit2d_cnt_pooling_a1 = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1851" *) 1'b1;
  assign unit2d_cnt_pooling_a2 = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1852" *) 2'b10;
  assign unit2d_cnt_pooling_a3 = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1853" *) 2'b11;
  assign unit2d_cnt_pooling_a4 = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1854" *) 3'b100;
  assign unit2d_cnt_pooling_a5 = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1855" *) 3'b101;
  assign unit2d_cnt_pooling_a6 = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1856" *) 3'b110;
  assign unit2d_cnt_pooling_a7 = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1857" *) 3'b111;
  assign _1239_ = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1879" *) 1'b1;
  assign _1240_ = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1888" *) 2'b10;
  assign _1241_ = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1897" *) 2'b11;
  assign _1242_ = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1906" *) 3'b100;
  assign _1243_ = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1915" *) 3'b101;
  assign _1244_ = unit2d_cnt_pooling + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1924" *) 3'b110;
  assign _1245_ = channel_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2111" *) 1'b1;
  assign _1246_ = line_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2126" *) 1'b1;
  assign _1247_ = bubble_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2140" *) 1'b1;
  assign _1248_ = last_out_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2185" *) 1'b1;
  assign _1249_ = one_width_bubble_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2280" *) 1'b1;
  assign _1250_ = unit2d_cnt_stride + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2302" *) 1'b1;
  assign rest_height_use = rest_height + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2327" *) reg2dp_pad_bottom_cfg;
  assign _1251_ = unit2d_vsize_cnt_0 + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2655" *) 1'b1;
  assign _1252_ = unit2d_vsize_cnt_1 + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2665" *) 1'b1;
  assign _1253_ = unit2d_vsize_cnt_2 + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2675" *) 1'b1;
  assign _1254_ = unit2d_vsize_cnt_3 + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2685" *) 1'b1;
  assign _1255_ = unit2d_vsize_cnt_4 + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2695" *) 1'b1;
  assign _1256_ = unit2d_vsize_cnt_5 + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2705" *) 1'b1;
  assign _1257_ = unit2d_vsize_cnt_6 + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2715" *) 1'b1;
  assign _1258_ = unit2d_vsize_cnt_7 + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2725" *) 1'b1;
  assign _1259_ = wr_sub_lbuf_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3423" *) 1'b1;
  assign _1260_ = sub_lbuf_dout_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3436" *) 1'b1;
  assign _0664_ = $signed(_0658_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0656_);
  assign _0744_ = $signed(_0738_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0736_);
  assign _0824_ = $signed(_0818_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0816_);
  assign _0904_ = $signed(_0898_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0896_);
  assign _0674_ = $signed(_0668_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0666_);
  assign _0754_ = $signed(_0748_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0746_);
  assign _0834_ = $signed(_0828_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0826_);
  assign _0914_ = $signed(_0908_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0906_);
  assign _0684_ = $signed(_0678_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0676_);
  assign _0764_ = $signed(_0758_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0756_);
  assign _0844_ = $signed(_0838_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0836_);
  assign _0924_ = $signed(_0918_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0916_);
  assign _0694_ = $signed(_0688_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0686_);
  assign _0774_ = $signed(_0768_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0766_);
  assign _0854_ = $signed(_0848_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0846_);
  assign _0934_ = $signed(_0928_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0926_);
  assign _0704_ = $signed(_0698_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0696_);
  assign _0784_ = $signed(_0778_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0776_);
  assign _0864_ = $signed(_0858_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0856_);
  assign _0944_ = $signed(_0938_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0936_);
  assign _0714_ = $signed(_0708_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0706_);
  assign _0794_ = $signed(_0788_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0786_);
  assign _0874_ = $signed(_0868_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0866_);
  assign _0954_ = $signed(_0948_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0946_);
  assign _0724_ = $signed(_0718_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0716_);
  assign _0804_ = $signed(_0798_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0796_);
  assign _0884_ = $signed(_0878_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0876_);
  assign _0964_ = $signed(_0958_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0956_);
  assign _0734_ = $signed(_0728_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0726_);
  assign _0814_ = $signed(_0808_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0806_);
  assign _0894_ = $signed(_0888_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0886_);
  assign _0974_ = $signed(_0968_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3557" *) $signed(_0966_);
  assign _0665_ = $signed(_0659_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0657_);
  assign _0745_ = $signed(_0739_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0737_);
  assign _0825_ = $signed(_0819_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0817_);
  assign _0905_ = $signed(_0899_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0897_);
  assign _0675_ = $signed(_0669_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0667_);
  assign _0755_ = $signed(_0749_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0747_);
  assign _0835_ = $signed(_0829_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0827_);
  assign _0915_ = $signed(_0909_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0907_);
  assign _0685_ = $signed(_0679_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0677_);
  assign _0765_ = $signed(_0759_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0757_);
  assign _0845_ = $signed(_0839_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0837_);
  assign _0925_ = $signed(_0919_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0917_);
  assign _0695_ = $signed(_0689_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0687_);
  assign _0775_ = $signed(_0769_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0767_);
  assign _0855_ = $signed(_0849_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0847_);
  assign _0935_ = $signed(_0929_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0927_);
  assign _0705_ = $signed(_0699_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0697_);
  assign _0785_ = $signed(_0779_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0777_);
  assign _0865_ = $signed(_0859_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0857_);
  assign _0945_ = $signed(_0939_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0937_);
  assign _0715_ = $signed(_0709_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0707_);
  assign _0795_ = $signed(_0789_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0787_);
  assign _0875_ = $signed(_0869_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0867_);
  assign _0955_ = $signed(_0949_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0947_);
  assign _0725_ = $signed(_0719_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0717_);
  assign _0805_ = $signed(_0799_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0797_);
  assign _0885_ = $signed(_0879_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0877_);
  assign _0965_ = $signed(_0959_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0957_);
  assign _0735_ = $signed(_0729_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0727_);
  assign _0815_ = $signed(_0809_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0807_);
  assign _0895_ = $signed(_0889_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0887_);
  assign _0975_ = $signed(_0969_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3558" *) $signed(_0967_);
  assign _0663_ = $signed(_0661_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0660_);
  assign _0743_ = $signed(_0741_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0740_);
  assign _0823_ = $signed(_0821_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0820_);
  assign _0903_ = $signed(_0901_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0900_);
  assign _0673_ = $signed(_0671_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0670_);
  assign _0753_ = $signed(_0751_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0750_);
  assign _0833_ = $signed(_0831_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0830_);
  assign _0913_ = $signed(_0911_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0910_);
  assign _0683_ = $signed(_0681_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0680_);
  assign _0763_ = $signed(_0761_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0760_);
  assign _0843_ = $signed(_0841_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0840_);
  assign _0923_ = $signed(_0921_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0920_);
  assign _0693_ = $signed(_0691_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0690_);
  assign _0773_ = $signed(_0771_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0770_);
  assign _0853_ = $signed(_0851_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0850_);
  assign _0933_ = $signed(_0931_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0930_);
  assign _0703_ = $signed(_0701_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0700_);
  assign _0783_ = $signed(_0781_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0780_);
  assign _0863_ = $signed(_0861_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0860_);
  assign _0943_ = $signed(_0941_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0940_);
  assign _0713_ = $signed(_0711_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0710_);
  assign _0793_ = $signed(_0791_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0790_);
  assign _0873_ = $signed(_0871_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0870_);
  assign _0953_ = $signed(_0951_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0950_);
  assign _0723_ = $signed(_0721_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0720_);
  assign _0803_ = $signed(_0801_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0800_);
  assign _0883_ = $signed(_0881_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0880_);
  assign _0963_ = $signed(_0961_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0960_);
  assign _0733_ = $signed(_0731_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0730_);
  assign _0813_ = $signed(_0811_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0810_);
  assign _0893_ = $signed(_0891_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0890_);
  assign _0973_ = $signed(_0971_) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3559" *) $signed(_0970_);
  assign _1261_ = unit2d_cnt_pooling_last + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5045" *) 1'b1;
  assign _1262_ = rd_line_out_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5813" *) 1'b1;
  assign _1263_ = rd_sub_lbuf_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5825" *) 1'b1;
  assign _1264_[2:0] = rd_comb_lbuf_cnt + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5838" *) 1'b1;
  assign kernel_width_cfg = reg2dp_kernel_width + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6288" *) 1'b1;
  assign data_16bit_0_ff = $signed(pout_mem_data_0[21:0]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6294" *) $signed(pad_value);
  assign data_16bit_1_ff = $signed(pout_mem_data_1[21:0]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6295" *) $signed(pad_value);
  assign data_16bit_2_ff = $signed(pout_mem_data_2[21:0]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6296" *) $signed(pad_value);
  assign data_16bit_3_ff = $signed(pout_mem_data_3[21:0]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6297" *) $signed(pad_value);
  assign data_8bit_0_ff = $signed(pout_mem_data_0[13:0]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6302" *) $signed(pad_value[13:0]);
  assign data_8bit_1_ff = $signed(pout_mem_data_0[27:14]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6303" *) $signed(pad_value[13:0]);
  assign data_8bit_2_ff = $signed(pout_mem_data_1[13:0]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6304" *) $signed(pad_value[13:0]);
  assign data_8bit_3_ff = $signed(pout_mem_data_1[27:14]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6305" *) $signed(pad_value[13:0]);
  assign data_8bit_4_ff = $signed(pout_mem_data_2[13:0]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6306" *) $signed(pad_value[13:0]);
  assign data_8bit_5_ff = $signed(pout_mem_data_2[27:14]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6307" *) $signed(pad_value[13:0]);
  assign data_8bit_6_ff = $signed(pout_mem_data_3[13:0]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6308" *) $signed(pad_value[13:0]);
  assign data_8bit_7_ff = $signed(pout_mem_data_3[27:14]) + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6309" *) $signed(pad_value[13:0]);
  assign i16_neg_add1_0 = data_hmult_16bit_0_ext[34:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6382" *) 1'b1;
  assign i16_neg_add1_1 = data_hmult_16bit_1_ext[34:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6383" *) 1'b1;
  assign i16_neg_add1_2 = data_hmult_16bit_2_ext[34:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6384" *) 1'b1;
  assign i16_neg_add1_3 = data_hmult_16bit_3_ext[34:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6385" *) 1'b1;
  assign _1265_ = data_hmult_16bit_0_ext[33:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6386" *) data_hmult_16bit_0_ext[15];
  assign _1266_ = data_hmult_16bit_1_ext[33:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6387" *) data_hmult_16bit_1_ext[15];
  assign _1267_ = data_hmult_16bit_2_ext[33:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6388" *) data_hmult_16bit_2_ext[15];
  assign _1268_ = data_hmult_16bit_3_ext[33:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6389" *) data_hmult_16bit_3_ext[15];
  assign i8_neg_add1_0_l = data_hmult_8bit_0_lsb_ext[26:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6603" *) 1'b1;
  assign i8_neg_add1_0_m = data_hmult_8bit_0_msb_ext[26:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6604" *) 1'b1;
  assign i8_neg_add1_1_l = data_hmult_8bit_1_lsb_ext[26:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6605" *) 1'b1;
  assign i8_neg_add1_1_m = data_hmult_8bit_1_msb_ext[26:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6606" *) 1'b1;
  assign i8_neg_add1_2_l = data_hmult_8bit_2_lsb_ext[26:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6607" *) 1'b1;
  assign i8_neg_add1_2_m = data_hmult_8bit_2_msb_ext[26:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6608" *) 1'b1;
  assign i8_neg_add1_3_l = data_hmult_8bit_3_lsb_ext[26:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6609" *) 1'b1;
  assign i8_neg_add1_3_m = data_hmult_8bit_3_msb_ext[26:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6610" *) 1'b1;
  assign _1269_ = data_hmult_8bit_0_lsb_ext[25:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6611" *) data_hmult_8bit_0_lsb_ext[15];
  assign _1270_ = data_hmult_8bit_0_msb_ext[25:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6612" *) data_hmult_8bit_0_msb_ext[15];
  assign _1271_ = data_hmult_8bit_1_lsb_ext[25:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6613" *) data_hmult_8bit_1_lsb_ext[15];
  assign _1272_ = data_hmult_8bit_1_msb_ext[25:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6614" *) data_hmult_8bit_1_msb_ext[15];
  assign _1273_ = data_hmult_8bit_2_lsb_ext[25:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6615" *) data_hmult_8bit_2_lsb_ext[15];
  assign _1274_ = data_hmult_8bit_2_msb_ext[25:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6616" *) data_hmult_8bit_2_msb_ext[15];
  assign _1275_ = data_hmult_8bit_3_lsb_ext[25:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6617" *) data_hmult_8bit_3_lsb_ext[15];
  assign _1276_ = data_hmult_8bit_3_msb_ext[25:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6618" *) data_hmult_8bit_3_msb_ext[15];
  assign i16_neg_vadd1_0 = data_vmult_16bit_0_ext[31:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7037" *) 1'b1;
  assign i16_neg_vadd1_1 = data_vmult_16bit_1_ext[31:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7038" *) 1'b1;
  assign i16_neg_vadd1_2 = data_vmult_16bit_2_ext[31:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7039" *) 1'b1;
  assign i16_neg_vadd1_3 = data_vmult_16bit_3_ext[31:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7040" *) 1'b1;
  assign _1277_ = data_vmult_16bit_0_ext[30:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7041" *) data_vmult_16bit_0_ext[15];
  assign _1278_ = data_vmult_16bit_1_ext[30:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7042" *) data_vmult_16bit_1_ext[15];
  assign _1279_ = data_vmult_16bit_2_ext[30:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7043" *) data_vmult_16bit_2_ext[15];
  assign _1280_ = data_vmult_16bit_3_ext[30:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7044" *) data_vmult_16bit_3_ext[15];
  assign i8_neg_vadd1_0_l = data_vmult_8bit_0_lsb_ext[23:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7258" *) 1'b1;
  assign i8_neg_vadd1_0_m = data_vmult_8bit_0_msb_ext[23:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7259" *) 1'b1;
  assign i8_neg_vadd1_1_l = data_vmult_8bit_1_lsb_ext[23:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7260" *) 1'b1;
  assign i8_neg_vadd1_1_m = data_vmult_8bit_1_msb_ext[23:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7261" *) 1'b1;
  assign i8_neg_vadd1_2_l = data_vmult_8bit_2_lsb_ext[23:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7262" *) 1'b1;
  assign i8_neg_vadd1_2_m = data_vmult_8bit_2_msb_ext[23:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7263" *) 1'b1;
  assign i8_neg_vadd1_3_l = data_vmult_8bit_3_lsb_ext[23:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7264" *) 1'b1;
  assign i8_neg_vadd1_3_m = data_vmult_8bit_3_msb_ext[23:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7265" *) 1'b1;
  assign _1281_ = data_vmult_8bit_0_lsb_ext[22:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7266" *) data_vmult_8bit_0_lsb_ext[15];
  assign _1282_ = data_vmult_8bit_0_msb_ext[22:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7267" *) data_vmult_8bit_0_msb_ext[15];
  assign _1283_ = data_vmult_8bit_1_lsb_ext[22:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7268" *) data_vmult_8bit_1_lsb_ext[15];
  assign _1284_ = data_vmult_8bit_1_msb_ext[22:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7269" *) data_vmult_8bit_1_msb_ext[15];
  assign _1285_ = data_vmult_8bit_2_lsb_ext[22:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7270" *) data_vmult_8bit_2_lsb_ext[15];
  assign _1286_ = data_vmult_8bit_2_msb_ext[22:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7271" *) data_vmult_8bit_2_msb_ext[15];
  assign _1287_ = data_vmult_8bit_3_lsb_ext[22:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7272" *) data_vmult_8bit_3_lsb_ext[15];
  assign _1288_ = data_vmult_8bit_3_msb_ext[22:16] + (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7273" *) data_vmult_8bit_3_msb_ext[15];
  assign pooling1d_prdy_use = one_width_norm_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1139" *) _2343_;
  assign one_width_norm_rdy = pooling1d_norm_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1140" *) _2344_;
  assign load_din = pooling1d_prdy_use & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1142" *) pooling1d_pvld;
  assign stripe_receive_done = load_din & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1143" *) data_c_end;
  assign wr_line_dat_done = _2011_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1168" *) stripe_receive_done;
  assign wr_surface_dat_done = wr_line_dat_done & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1181" *) last_line_in;
  assign wr_subcube_dat_done = _2012_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1201" *) wr_surface_dat_done;
  assign wr_total_cube_done = _2013_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1213" *) wr_subcube_dat_done;
  assign last_splitw = _2013_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1217" *) splitw_enable;
  assign first_splitw = _2014_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1218" *) splitw_enable;
  assign middle_surface_trig = wr_surface_dat_done & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1301" *) _2345_;
  assign stride_end = wr_line_dat_done & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1302" *) _2015_;
  assign small_active = _2346_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1440" *) _2339_;
  assign _1289_ = wr_subcube_dat_done & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2055" *) need_flush;
  assign _1290_ = _1289_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2055" *) is_one_width_in;
  assign _1291_ = wr_surface_dat_done & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2065" *) need_bubble;
  assign _1292_ = _1291_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2065" *) is_one_width_in;
  assign _1293_ = _1289_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2076" *) _2347_;
  assign _1294_ = subend_need_flush_flg & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2076" *) one_width_bubble_end;
  assign _1295_ = _1291_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2078" *) _2347_;
  assign _1296_ = surfend_need_bubble_flg & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2078" *) one_width_bubble_end;
  assign last_c = _2214_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2117" *) one_width_norm_rdy;
  assign line_end = _2215_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2131" *) last_c;
  assign bubble_en_end = _2216_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2145" *) line_end;
  assign _1297_ = need_bubble & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) bubble_en_end;
  assign _1298_ = _1297_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) _2348_;
  assign _1299_ = _1298_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) _2340_;
  assign _1300_ = _2349_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) need_flush;
  assign _1301_ = _1300_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) wr_surface_dat_done;
  assign _1302_ = _1301_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) _2350_;
  assign _1303_ = _2217_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2182" *) need_bubble;
  assign _1304_ = _2349_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2182" *) _2218_;
  assign _1305_ = _2622_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2237" *) wr_line_dat_done;
  assign last_out_done = _1305_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2237" *) last_out_en;
  assign _1306_ = wr_line_dat_done & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2265" *) is_one_width_in;
  assign one_width_bubble_end = _2223_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2285" *) pooling1d_norm_rdy;
  assign pooling_2d_rdy = wr_line_dat_done & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2287" *) _2224_;
  assign init_unit2d_set[0] = init_cnt & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2331" *) _2289_;
  assign _1307_ = stride_end & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2332" *) stride_trig_end;
  assign unit2d_set_trig[0] = _1307_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2332" *) _2351_;
  assign _1308_ = pooling_2d_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2334" *) _2225_;
  assign init_unit2d_set[1] = init_cnt & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2347" *) _2290_;
  assign _1309_ = stride_end & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2348" *) _2226_;
  assign _1310_ = _1309_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2348" *) _2352_;
  assign unit2d_set_trig[1] = _1310_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2348" *) _2351_;
  assign _1311_ = pooling_2d_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2350" *) _2227_;
  assign init_unit2d_set[2] = init_cnt & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2363" *) _2291_;
  assign _1312_ = stride_end & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2364" *) _2228_;
  assign _1313_ = _1312_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2364" *) _2352_;
  assign unit2d_set_trig[2] = _1313_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2364" *) _2351_;
  assign _1314_ = pooling_2d_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2366" *) _2229_;
  assign init_unit2d_set[3] = init_cnt & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2379" *) _2292_;
  assign _1315_ = stride_end & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2380" *) _2230_;
  assign _1316_ = _1315_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2380" *) _2352_;
  assign unit2d_set_trig[3] = _1316_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2380" *) _2351_;
  assign _1317_ = pooling_2d_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2382" *) _2231_;
  assign init_unit2d_set[4] = init_cnt & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2395" *) _2293_;
  assign _1318_ = stride_end & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2396" *) _2232_;
  assign _1319_ = _1318_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2396" *) _2352_;
  assign unit2d_set_trig[4] = _1319_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2396" *) _2351_;
  assign _1320_ = pooling_2d_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2398" *) _2233_;
  assign init_unit2d_set[5] = init_cnt & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2411" *) _2294_;
  assign _1321_ = stride_end & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2412" *) _2234_;
  assign _1322_ = _1321_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2412" *) _2352_;
  assign unit2d_set_trig[5] = _1322_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2412" *) _2351_;
  assign _1323_ = pooling_2d_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2414" *) _2235_;
  assign init_unit2d_set[6] = init_cnt & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2427" *) _2295_;
  assign _1324_ = stride_end & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2428" *) _2236_;
  assign _1325_ = _1324_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2428" *) _2352_;
  assign unit2d_set_trig[6] = _1325_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2428" *) _2351_;
  assign _1326_ = pooling_2d_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2430" *) _2237_;
  assign init_unit2d_set[7] = init_cnt & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2443" *) _2296_;
  assign _1327_ = stride_end & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2444" *) _2238_;
  assign _1328_ = _1327_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2444" *) _2352_;
  assign unit2d_set_trig[7] = _1328_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2444" *) _2351_;
  assign _1329_ = pooling_2d_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2446" *) _2239_;
  assign _1330_ = unit2d_en[0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2654" *) wr_line_dat_done;
  assign _1331_ = unit2d_en[1] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2664" *) wr_line_dat_done;
  assign _1332_ = unit2d_en[2] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2674" *) wr_line_dat_done;
  assign _1333_ = unit2d_en[3] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2684" *) wr_line_dat_done;
  assign _1334_ = unit2d_en[4] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2694" *) wr_line_dat_done;
  assign _1335_ = unit2d_en[5] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2704" *) wr_line_dat_done;
  assign _1336_ = unit2d_en[6] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2714" *) wr_line_dat_done;
  assign _1337_ = unit2d_en[7] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2724" *) wr_line_dat_done;
  assign _1338_ = unit2d_en[0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3327" *) load_din;
  assign _1339_ = _1338_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3327" *) _2240_;
  assign mem_re1[0] = _1339_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3327" *) mem_re1_sel;
  assign _1340_ = _1338_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3328" *) _2241_;
  assign mem_re1[1] = _1340_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3328" *) mem_re1_sel;
  assign _1341_ = _1338_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3329" *) _2242_;
  assign mem_re1[2] = _1341_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3329" *) mem_re1_sel;
  assign _1342_ = _1338_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3330" *) _2243_;
  assign mem_re1[3] = _1342_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3330" *) mem_re1_sel;
  assign _1343_ = _1338_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3331" *) _2244_;
  assign mem_re1[4] = _1343_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3331" *) mem_re1_sel;
  assign _1344_ = _1338_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3332" *) _2245_;
  assign mem_re1[5] = _1344_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3332" *) mem_re1_sel;
  assign _1345_ = _1338_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3333" *) _2246_;
  assign mem_re1[6] = _1345_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3333" *) mem_re1_sel;
  assign _1346_ = _1338_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3334" *) _2247_;
  assign mem_re1[7] = _1346_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3334" *) mem_re1_sel;
  assign mem_re1_1st[7] = unit2d_mem_1strd[0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3335" *) mem_re1_sel;
  assign mem_re2[0] = _1339_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3346" *) mem_re2_sel;
  assign mem_re2[1] = _1340_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3347" *) mem_re2_sel;
  assign mem_re2[2] = _1341_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3348" *) mem_re2_sel;
  assign mem_re2[3] = _1342_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3349" *) mem_re2_sel;
  assign _1347_ = unit2d_en[1] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3350" *) load_din;
  assign _1348_ = _1347_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3350" *) _2240_;
  assign mem_re2[4] = _1348_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3350" *) mem_re2_sel;
  assign _1349_ = _1347_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3351" *) _2241_;
  assign mem_re2[5] = _1349_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3351" *) mem_re2_sel;
  assign _1350_ = _1347_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3352" *) _2242_;
  assign mem_re2[6] = _1350_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3352" *) mem_re2_sel;
  assign _1351_ = _1347_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3353" *) _2243_;
  assign mem_re2[7] = _1351_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3353" *) mem_re2_sel;
  assign mem_re2_1st[3] = unit2d_mem_1strd[0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3354" *) mem_re2_sel;
  assign mem_re2_1st[7] = unit2d_mem_1strd[1] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3358" *) mem_re2_sel;
  assign mem_re3[0] = _1339_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3363" *) mem_re3_sel;
  assign mem_re3[1] = _1340_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3364" *) mem_re3_sel;
  assign mem_re3[2] = _1348_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3365" *) mem_re3_sel;
  assign mem_re3[3] = _1349_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3366" *) mem_re3_sel;
  assign _1352_ = unit2d_en[2] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3367" *) load_din;
  assign _1353_ = _1352_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3367" *) _2240_;
  assign mem_re3[4] = _1353_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3367" *) mem_re3_sel;
  assign _1354_ = _1352_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3368" *) _2241_;
  assign mem_re3[5] = _1354_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3368" *) mem_re3_sel;
  assign _1355_ = unit2d_en[3] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3369" *) load_din;
  assign _1356_ = _1355_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3369" *) _2240_;
  assign mem_re3[6] = _1356_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3369" *) mem_re3_sel;
  assign _1357_ = _1355_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3370" *) _2241_;
  assign mem_re3[7] = _1357_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3370" *) mem_re3_sel;
  assign mem_re3_1st[1] = unit2d_mem_1strd[0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3371" *) mem_re3_sel;
  assign mem_re3_1st[3] = unit2d_mem_1strd[1] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3373" *) mem_re3_sel;
  assign mem_re3_1st[5] = unit2d_mem_1strd[2] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3375" *) mem_re3_sel;
  assign mem_re3_1st[7] = unit2d_mem_1strd[3] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3377" *) mem_re3_sel;
  assign mem_re4[0] = _1339_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3380" *) mem_re4_sel;
  assign mem_re4[1] = _1348_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3381" *) mem_re4_sel;
  assign mem_re4[2] = _1353_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3382" *) mem_re4_sel;
  assign mem_re4[3] = _1356_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3383" *) mem_re4_sel;
  assign _1358_ = unit2d_en[4] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3384" *) load_din;
  assign _1359_ = _1358_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3384" *) _2240_;
  assign mem_re4[4] = _1359_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3384" *) mem_re4_sel;
  assign _1360_ = unit2d_en[5] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3385" *) load_din;
  assign _1361_ = _1360_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3385" *) _2240_;
  assign mem_re4[5] = _1361_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3385" *) mem_re4_sel;
  assign _1362_ = unit2d_en[6] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3386" *) load_din;
  assign _1363_ = _1362_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3386" *) _2240_;
  assign mem_re4[6] = _1363_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3386" *) mem_re4_sel;
  assign _1364_ = unit2d_en[7] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3387" *) load_din;
  assign _1365_ = _1364_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3387" *) _2240_;
  assign mem_re4[7] = _1365_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3387" *) mem_re4_sel;
  assign mem_re4_1st[0] = unit2d_mem_1strd[0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3388" *) mem_re4_sel;
  assign mem_re4_1st[1] = unit2d_mem_1strd[1] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3389" *) mem_re4_sel;
  assign mem_re4_1st[2] = unit2d_mem_1strd[2] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3390" *) mem_re4_sel;
  assign mem_re4_1st[3] = unit2d_mem_1strd[3] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3391" *) mem_re4_sel;
  assign mem_re4_1st[4] = unit2d_mem_1strd[4] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3392" *) mem_re4_sel;
  assign mem_re4_1st[5] = unit2d_mem_1strd[5] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3393" *) mem_re4_sel;
  assign mem_re4_1st[6] = unit2d_mem_1strd[6] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3394" *) mem_re4_sel;
  assign mem_re4_1st[7] = unit2d_mem_1strd[7] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3395" *) mem_re4_sel;
  assign last_sub_lbuf_done = _2250_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3426" *) sub_lbuf_dout_done;
  assign _1366_ = cur_datin_disable & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3435" *) one_width_norm_rdy;
  assign sub_lbuf_dout_done = _2251_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3440" *) _2262_;
  assign _1367_ = _0403_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[0];
  assign _1368_ = _0467_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[0];
  assign _1369_ = _0531_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[0];
  assign _1370_ = _0595_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[0];
  assign _1371_ = _0411_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[1];
  assign _1372_ = _0475_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[1];
  assign _1373_ = _0539_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[1];
  assign _1374_ = _0603_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[1];
  assign _1375_ = _0419_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[2];
  assign _1376_ = _0483_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[2];
  assign _1377_ = _0547_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[2];
  assign _1378_ = _0611_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[2];
  assign _1379_ = _0427_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[3];
  assign _1380_ = _0491_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[3];
  assign _1381_ = _0555_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[3];
  assign _1382_ = _0619_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[3];
  assign _1383_ = _0435_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[4];
  assign _1384_ = _0499_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[4];
  assign _1385_ = _0563_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[4];
  assign _1386_ = _0627_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[4];
  assign _1387_ = _0443_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[5];
  assign _1388_ = _0507_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[5];
  assign _1389_ = _0571_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[5];
  assign _1390_ = _0635_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[5];
  assign _1391_ = _0451_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[6];
  assign _1392_ = _0515_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[6];
  assign _1393_ = _0579_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[6];
  assign _1394_ = _0643_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[6];
  assign _1395_ = _0459_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[7];
  assign _1396_ = _0523_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[7];
  assign _1397_ = _0587_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[7];
  assign _1398_ = _0651_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) mem_data_valid[7];
  assign _1399_ = _0405_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[0];
  assign _1400_ = _0469_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[0];
  assign _1401_ = _0533_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[0];
  assign _1402_ = _0597_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[0];
  assign _1403_ = _0413_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[1];
  assign _1404_ = _0477_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[1];
  assign _1405_ = _0541_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[1];
  assign _1406_ = _0605_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[1];
  assign _1407_ = _0421_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[2];
  assign _1408_ = _0485_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[2];
  assign _1409_ = _0549_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[2];
  assign _1410_ = _0613_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[2];
  assign _1411_ = _0429_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[3];
  assign _1412_ = _0493_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[3];
  assign _1413_ = _0557_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[3];
  assign _1414_ = _0621_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[3];
  assign _1415_ = _0437_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[4];
  assign _1416_ = _0501_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[4];
  assign _1417_ = _0565_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[4];
  assign _1418_ = _0629_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[4];
  assign _1419_ = _0445_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[5];
  assign _1420_ = _0509_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[5];
  assign _1421_ = _0573_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[5];
  assign _1422_ = _0637_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[5];
  assign _1423_ = _0453_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[6];
  assign _1424_ = _0517_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[6];
  assign _1425_ = _0581_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[6];
  assign _1426_ = _0645_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[6];
  assign _1427_ = _0461_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[7];
  assign _1428_ = _0525_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[7];
  assign _1429_ = _0589_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[7];
  assign _1430_ = _0653_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) mem_data_valid[7];
  assign _1431_ = _0401_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[0];
  assign _1432_ = _0465_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[0];
  assign _1433_ = _0529_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[0];
  assign _1434_ = _0593_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[0];
  assign _1435_ = _0409_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[1];
  assign _1436_ = _0473_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[1];
  assign _1437_ = _0537_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[1];
  assign _1438_ = _0601_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[1];
  assign _1439_ = _0417_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[2];
  assign _1440_ = _0481_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[2];
  assign _1441_ = _0545_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[2];
  assign _1442_ = _0609_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[2];
  assign _1443_ = _0425_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[3];
  assign _1444_ = _0489_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[3];
  assign _1445_ = _0553_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[3];
  assign _1446_ = _0617_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[3];
  assign _1447_ = _0433_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[4];
  assign _1448_ = _0497_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[4];
  assign _1449_ = _0561_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[4];
  assign _1450_ = _0625_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[4];
  assign _1451_ = _0441_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[5];
  assign _1452_ = _0505_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[5];
  assign _1453_ = _0569_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[5];
  assign _1454_ = _0633_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[5];
  assign _1455_ = _0449_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[6];
  assign _1456_ = _0513_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[6];
  assign _1457_ = _0577_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[6];
  assign _1458_ = _0641_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[6];
  assign _1459_ = _0457_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[7];
  assign _1460_ = _0521_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[7];
  assign _1461_ = _0585_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[7];
  assign _1462_ = _0649_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) mem_data_valid[7];
  assign _1463_ = _2353_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2354_;
  assign _1464_ = _2355_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2356_;
  assign _1465_ = _2357_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2358_;
  assign _1466_ = _2359_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2360_;
  assign _1467_ = _2353_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2361_;
  assign _1468_ = _2355_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2362_;
  assign _1469_ = _2357_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2363_;
  assign _1470_ = _2359_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2364_;
  assign _1471_ = _2353_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2365_;
  assign _1472_ = _2355_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2366_;
  assign _1473_ = _2357_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2367_;
  assign _1474_ = _2359_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2368_;
  assign _1475_ = _2353_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2369_;
  assign _1476_ = _2355_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2370_;
  assign _1477_ = _2357_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2371_;
  assign _1478_ = _2359_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2372_;
  assign _1479_ = _2353_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2373_;
  assign _1480_ = _2355_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2374_;
  assign _1481_ = _2357_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2375_;
  assign _1482_ = _2359_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2376_;
  assign _1483_ = _2353_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2377_;
  assign _1484_ = _2355_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2378_;
  assign _1485_ = _2357_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2379_;
  assign _1486_ = _2359_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2380_;
  assign _1487_ = _2353_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2381_;
  assign _1488_ = _2355_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2382_;
  assign _1489_ = _2357_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2383_;
  assign _1490_ = _2359_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2384_;
  assign _1491_ = _2353_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2385_;
  assign _1492_ = _2355_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2386_;
  assign _1493_ = _2357_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2387_;
  assign _1494_ = _2359_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _2388_;
  assign _1495_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0005_[15];
  assign _1496_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0105_[15];
  assign _1497_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0205_[15];
  assign _1498_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0305_[15];
  assign _1499_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0018_[15];
  assign _1500_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0118_[15];
  assign _1501_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0218_[15];
  assign _1502_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0318_[15];
  assign _1503_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0030_[15];
  assign _1504_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0130_[15];
  assign _1505_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0230_[15];
  assign _1506_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0330_[15];
  assign _1507_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0042_[15];
  assign _1508_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0142_[15];
  assign _1509_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0242_[15];
  assign _1510_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0342_[15];
  assign _1511_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0054_[15];
  assign _1512_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0154_[15];
  assign _1513_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0254_[15];
  assign _1514_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0354_[15];
  assign _1515_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0066_[15];
  assign _1516_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0166_[15];
  assign _1517_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0266_[15];
  assign _1518_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0366_[15];
  assign _1519_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0078_[15];
  assign _1520_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0178_[15];
  assign _1521_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0278_[15];
  assign _1522_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0378_[15];
  assign _1523_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0090_[15];
  assign _1524_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0190_[15];
  assign _1525_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0290_[15];
  assign _1526_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0390_[15];
  assign _1527_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2354_;
  assign _1528_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2356_;
  assign _1529_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2358_;
  assign _1530_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2360_;
  assign _1531_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2361_;
  assign _1532_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2362_;
  assign _1533_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2363_;
  assign _1534_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2364_;
  assign _1535_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2365_;
  assign _1536_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2366_;
  assign _1537_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2367_;
  assign _1538_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2368_;
  assign _1539_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2369_;
  assign _1540_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2370_;
  assign _1541_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2371_;
  assign _1542_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2372_;
  assign _1543_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2373_;
  assign _1544_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2374_;
  assign _1545_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2375_;
  assign _1546_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2376_;
  assign _1547_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2377_;
  assign _1548_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2378_;
  assign _1549_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2379_;
  assign _1550_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2380_;
  assign _1551_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2381_;
  assign _1552_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2382_;
  assign _1553_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2383_;
  assign _1554_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2384_;
  assign _1555_ = _0004_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2385_;
  assign _1556_ = _0104_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _2386_;
  assign _1559_ = _0011_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[0];
  assign _1560_ = _0111_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[0];
  assign _1561_ = _0211_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[0];
  assign _1562_ = _0311_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[0];
  assign _1563_ = _0023_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[1];
  assign _1564_ = _0123_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[1];
  assign _1565_ = _0223_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[1];
  assign _1566_ = _0323_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[1];
  assign _1567_ = _0035_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[2];
  assign _1568_ = _0135_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[2];
  assign _1569_ = _0235_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[2];
  assign _1570_ = _0335_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[2];
  assign _1571_ = _0047_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[3];
  assign _1572_ = _0147_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[3];
  assign _1573_ = _0247_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[3];
  assign _1574_ = _0347_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[3];
  assign _1575_ = _0059_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[4];
  assign _1576_ = _0159_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[4];
  assign _1577_ = _0259_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[4];
  assign _1578_ = _0359_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[4];
  assign _1579_ = _0071_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[5];
  assign _1580_ = _0171_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[5];
  assign _1581_ = _0271_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[5];
  assign _1582_ = _0371_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[5];
  assign _1583_ = _0083_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[6];
  assign _1584_ = _0183_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[6];
  assign _1585_ = _0283_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[6];
  assign _1586_ = _0383_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[6];
  assign _1587_ = _0095_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[7];
  assign _1588_ = _0195_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[7];
  assign _1589_ = _0295_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[7];
  assign _1590_ = _0395_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) mem_data_valid[7];
  assign _1591_ = _0013_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[0];
  assign _1592_ = _0113_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[0];
  assign _1593_ = _0213_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[0];
  assign _1594_ = _0313_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[0];
  assign _1595_ = _0025_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[1];
  assign _1596_ = _0125_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[1];
  assign _1597_ = _0225_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[1];
  assign _1598_ = _0325_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[1];
  assign _1599_ = _0037_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[2];
  assign _1600_ = _0137_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[2];
  assign _1601_ = _0237_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[2];
  assign _1602_ = _0337_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[2];
  assign _1603_ = _0049_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[3];
  assign _1604_ = _0149_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[3];
  assign _1605_ = _0249_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[3];
  assign _1606_ = _0349_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[3];
  assign _1607_ = _0061_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[4];
  assign _1608_ = _0161_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[4];
  assign _1609_ = _0261_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[4];
  assign _1610_ = _0361_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[4];
  assign _1611_ = _0073_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[5];
  assign _1612_ = _0173_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[5];
  assign _1613_ = _0273_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[5];
  assign _1614_ = _0373_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[5];
  assign _1615_ = _0085_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[6];
  assign _1616_ = _0185_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[6];
  assign _1617_ = _0285_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[6];
  assign _1618_ = _0385_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[6];
  assign _1619_ = _0097_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[7];
  assign _1620_ = _0197_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[7];
  assign _1621_ = _0297_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[7];
  assign _1622_ = _0397_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) mem_data_valid[7];
  assign _1623_ = _0009_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[0];
  assign _1624_ = _0109_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[0];
  assign _1625_ = _0209_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[0];
  assign _1626_ = _0309_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[0];
  assign _1627_ = _0021_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[1];
  assign _1628_ = _0121_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[1];
  assign _1629_ = _0221_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[1];
  assign _1630_ = _0321_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[1];
  assign _1631_ = _0033_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[2];
  assign _1632_ = _0133_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[2];
  assign _1633_ = _0233_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[2];
  assign _1634_ = _0333_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[2];
  assign _1635_ = _0045_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[3];
  assign _1636_ = _0145_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[3];
  assign _1637_ = _0245_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[3];
  assign _1638_ = _0345_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[3];
  assign _1639_ = _0057_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[4];
  assign _1640_ = _0157_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[4];
  assign _1641_ = _0257_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[4];
  assign _1642_ = _0357_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[4];
  assign _1643_ = _0069_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[5];
  assign _1644_ = _0169_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[5];
  assign _1645_ = _0269_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[5];
  assign _1646_ = _0369_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[5];
  assign _1647_ = _0081_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[6];
  assign _1648_ = _0181_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[6];
  assign _1649_ = _0281_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[6];
  assign _1650_ = _0381_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[6];
  assign _1651_ = _0093_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[7];
  assign _1652_ = _0193_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[7];
  assign _1653_ = _0293_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[7];
  assign _1654_ = _0393_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) mem_data_valid[7];
  assign _1557_ = _0204_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _2387_;
  assign _1558_ = _0304_[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _2388_;
  assign _1655_ = reg2dp_int8_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) mem_data_valid[0];
  assign _1656_ = reg2dp_int8_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) mem_data_valid[1];
  assign _1657_ = reg2dp_int8_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) mem_data_valid[2];
  assign _1658_ = reg2dp_int8_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) mem_data_valid[3];
  assign _1659_ = reg2dp_int8_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) mem_data_valid[4];
  assign _1660_ = reg2dp_int8_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) mem_data_valid[5];
  assign _1661_ = reg2dp_int8_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) mem_data_valid[6];
  assign _1662_ = reg2dp_int8_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) mem_data_valid[7];
  assign _1663_ = reg2dp_int16_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) mem_data_valid[0];
  assign _1664_ = reg2dp_int16_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) mem_data_valid[1];
  assign _1665_ = reg2dp_int16_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) mem_data_valid[2];
  assign _1666_ = reg2dp_int16_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) mem_data_valid[3];
  assign _1667_ = reg2dp_int16_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) mem_data_valid[4];
  assign _1668_ = reg2dp_int16_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) mem_data_valid[5];
  assign _1669_ = reg2dp_int16_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) mem_data_valid[6];
  assign _1670_ = reg2dp_int16_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) mem_data_valid[7];
  assign _0977_[0] = _2980_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3586" *) _3074_;
  assign _0978_[0] = _2981_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) _3075_;
  assign _0983_[0] = _2982_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) _3076_;
  assign _0986_[0] = _2983_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) _3077_;
  assign _0989_[0] = _2984_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) _3078_;
  assign _0992_[0] = _2985_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) _3079_;
  assign _0995_[0] = _2986_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) _3080_;
  assign _0998_[0] = _2987_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) _3081_;
  assign _1001_[0] = _2988_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) _3082_;
  assign _0977_[1] = _2989_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3588" *) _3083_;
  assign _0978_[1] = _2990_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) _3084_;
  assign _0983_[1] = _2991_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) _3085_;
  assign _0986_[1] = _2992_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) _3086_;
  assign _0989_[1] = _2993_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) _3087_;
  assign _0992_[1] = _2994_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) _3088_;
  assign _0995_[1] = _2995_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) _3089_;
  assign _0998_[1] = _2996_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) _3090_;
  assign _1001_[1] = _2997_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) _3091_;
  assign _0977_[2] = _2998_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3590" *) _3092_;
  assign _0978_[2] = _2999_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) _3093_;
  assign _0983_[2] = _3000_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) _3094_;
  assign _0986_[2] = _3001_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) _3095_;
  assign _0989_[2] = _3002_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) _3096_;
  assign _0992_[2] = _3003_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) _3097_;
  assign _0995_[2] = _3004_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) _3098_;
  assign _0998_[2] = _3005_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) _3099_;
  assign _1001_[2] = _3006_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) _3100_;
  assign _0977_[3] = _3007_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3592" *) _3101_;
  assign _0978_[3] = _3008_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) _3102_;
  assign _0983_[3] = _3009_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) _3103_;
  assign _0986_[3] = _3010_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) _3104_;
  assign _0989_[3] = _3011_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) _3105_;
  assign _0992_[3] = _3012_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) _3106_;
  assign _0995_[3] = _3013_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) _3107_;
  assign _0998_[3] = _3014_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) _3108_;
  assign _1001_[3] = _3015_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) _3109_;
  assign _1671_ = _2390_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) reg2dp_fp16_en;
  assign _1672_ = _2391_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) reg2dp_fp16_en;
  assign _1673_ = _2392_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) reg2dp_fp16_en;
  assign _1674_ = _2393_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) reg2dp_fp16_en;
  assign _1675_ = _2394_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) reg2dp_fp16_en;
  assign _1676_ = _2395_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) reg2dp_fp16_en;
  assign _1677_ = _2396_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) reg2dp_fp16_en;
  assign _1678_ = _2397_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) reg2dp_fp16_en;
  assign _1679_ = _2398_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) reg2dp_fp16_en;
  assign _1680_ = _2399_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) reg2dp_fp16_en;
  assign _1681_ = _2400_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) reg2dp_fp16_en;
  assign _1682_ = _2401_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) reg2dp_fp16_en;
  assign _1683_ = _2402_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) reg2dp_fp16_en;
  assign _1684_ = _2403_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) reg2dp_fp16_en;
  assign _1685_ = _2404_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) reg2dp_fp16_en;
  assign _1686_ = _2405_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) reg2dp_fp16_en;
  assign _1687_ = _2406_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) reg2dp_fp16_en;
  assign _1688_ = _2407_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) reg2dp_fp16_en;
  assign _1689_ = _2408_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) reg2dp_fp16_en;
  assign _1690_ = _2409_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) reg2dp_fp16_en;
  assign _1691_ = _2410_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) reg2dp_fp16_en;
  assign _1692_ = _2411_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) reg2dp_fp16_en;
  assign _1693_ = _2412_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) reg2dp_fp16_en;
  assign _1694_ = _2413_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) reg2dp_fp16_en;
  assign _1695_ = _2414_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) reg2dp_fp16_en;
  assign _1696_ = _2415_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) reg2dp_fp16_en;
  assign _1697_ = _2416_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) reg2dp_fp16_en;
  assign _1698_ = _2417_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) reg2dp_fp16_en;
  assign _1699_ = _2418_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) reg2dp_fp16_en;
  assign _1700_ = _2419_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) reg2dp_fp16_en;
  assign _1701_ = _2420_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) reg2dp_fp16_en;
  assign _1702_ = _2421_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) reg2dp_fp16_en;
  assign _1703_ = flush_read_en_d & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3621" *) wr_data_stage0_prdy;
  assign _1704_ = flush_read_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4148" *) one_width_norm_rdy;
  assign load_din_all = pooling1d_norm_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4334" *) pooling1d_vld_rebuild;
  assign load_wr_stage1_all = wr_data_stage0_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4349" *) wr_data_stage0_prdy;
  assign _1705_ = load_wr_stage1_all & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4351" *) _2424_;
  assign load_wr_stage1 = _1705_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4351" *) _2425_;
  assign load_wr_stage2_all = wr_data_stage1_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4363" *) wr_data_stage1_prdy;
  assign _1706_ = load_wr_stage2_all & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4364" *) _2426_;
  assign load_wr_stage2 = _1706_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4364" *) _2427_;
  assign _1707_ = wr_data_stage1_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4370" *) _2428_;
  assign load_wr_stage3_all = wr_data_stage2_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4376" *) pout_data_stage0_prdy;
  assign _1708_ = load_wr_stage3_all & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4377" *) _2429_;
  assign load_wr_stage3 = _1708_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4377" *) _2430_;
  assign fp16_mean_pool_cfg = fp16_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4556" *) average_pooling_en;
  assign _1709_ = int_mem_we & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4566" *) { load_wr_stage3, load_wr_stage3, load_wr_stage3, load_wr_stage3, load_wr_stage3, load_wr_stage3, load_wr_stage3, load_wr_stage3 };
  assign _1710_ = line_end & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5041" *) cur_datin_disable;
  assign _1711_ = wr_line_dat_done & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5041" *) last_out_en;
  assign _1712_ = _2679_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5041" *) one_width_norm_rdy;
  assign flush_read_en = _2680_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5052" *) one_width_norm_rdy;
  assign unit2d_en_last[0] = flush_read_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5053" *) _2253_;
  assign unit2d_en_last[1] = flush_read_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5054" *) _2254_;
  assign unit2d_en_last[2] = flush_read_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5055" *) _2255_;
  assign unit2d_en_last[3] = flush_read_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5056" *) _2256_;
  assign unit2d_en_last[4] = flush_read_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5057" *) _2257_;
  assign unit2d_en_last[5] = flush_read_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5058" *) _2258_;
  assign unit2d_en_last[6] = flush_read_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5059" *) _2259_;
  assign unit2d_en_last[7] = flush_read_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5060" *) _2260_;
  assign _1713_ = unit2d_en_last[0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5061" *) _2240_;
  assign mem_re2_last[0] = _1713_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5061" *) mem_re2_sel_last;
  assign _1714_ = unit2d_en_last[0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5062" *) _2241_;
  assign mem_re2_last[1] = _1714_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5062" *) mem_re2_sel_last;
  assign _1715_ = unit2d_en_last[0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5063" *) _2242_;
  assign mem_re2_last[2] = _1715_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5063" *) mem_re2_sel_last;
  assign _1716_ = unit2d_en_last[0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5064" *) _2243_;
  assign mem_re2_last[3] = _1716_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5064" *) mem_re2_sel_last;
  assign _1717_ = unit2d_en_last[1] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5065" *) _2240_;
  assign mem_re2_last[4] = _1717_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5065" *) mem_re2_sel_last;
  assign _1718_ = unit2d_en_last[1] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5066" *) _2241_;
  assign mem_re2_last[5] = _1718_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5066" *) mem_re2_sel_last;
  assign _1719_ = unit2d_en_last[1] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5067" *) _2242_;
  assign mem_re2_last[6] = _1719_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5067" *) mem_re2_sel_last;
  assign _1720_ = unit2d_en_last[1] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5068" *) _2243_;
  assign mem_re2_last[7] = _1720_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5068" *) mem_re2_sel_last;
  assign mem_re3_last[0] = _1713_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5069" *) mem_re3_sel_last;
  assign mem_re3_last[1] = _1714_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5070" *) mem_re3_sel_last;
  assign mem_re3_last[2] = _1717_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5071" *) mem_re3_sel_last;
  assign mem_re3_last[3] = _1718_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5072" *) mem_re3_sel_last;
  assign _1721_ = unit2d_en_last[2] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5073" *) _2240_;
  assign mem_re3_last[4] = _1721_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5073" *) mem_re3_sel_last;
  assign _1722_ = unit2d_en_last[2] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5074" *) _2241_;
  assign mem_re3_last[5] = _1722_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5074" *) mem_re3_sel_last;
  assign _1723_ = unit2d_en_last[3] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5075" *) _2240_;
  assign mem_re3_last[6] = _1723_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5075" *) mem_re3_sel_last;
  assign _1724_ = unit2d_en_last[3] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5076" *) _2241_;
  assign mem_re3_last[7] = _1724_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5076" *) mem_re3_sel_last;
  assign mem_re4_last[0] = _1713_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5077" *) mem_re4_sel_last;
  assign mem_re4_last[1] = _1717_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5078" *) mem_re4_sel_last;
  assign mem_re4_last[2] = _1721_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5079" *) mem_re4_sel_last;
  assign mem_re4_last[3] = _1723_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5080" *) mem_re4_sel_last;
  assign _1725_ = unit2d_en_last[4] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5081" *) _2240_;
  assign mem_re4_last[4] = _1725_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5081" *) mem_re4_sel_last;
  assign _1726_ = unit2d_en_last[5] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5082" *) _2240_;
  assign mem_re4_last[5] = _1726_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5082" *) mem_re4_sel_last;
  assign _1727_ = unit2d_en_last[6] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5083" *) _2240_;
  assign mem_re4_last[6] = _1727_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5083" *) mem_re4_sel_last;
  assign _1728_ = unit2d_en_last[7] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5084" *) _2240_;
  assign mem_re4_last[7] = _1728_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5084" *) mem_re4_sel_last;
  assign _1729_ = load_din & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5090" *) _3111_;
  assign _1730_ = cur_datin_disable_d & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5395" *) wr_data_stage0_prdy;
  assign _1731_ = load_wr_stage1 & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5456" *) _3112_;
  assign _1732_ = cur_datin_disable_2d & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5764" *) wr_data_stage1_prdy;
  assign _1733_ = _2682_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5764" *) mem_re_last_2d[0];
  assign _1734_ = _1733_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5764" *) _2265_;
  assign pout_mem_data_sel_1_last[0] = _1734_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5764" *) mem_re2_sel;
  assign _1735_ = _2682_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5765" *) mem_re_last_2d[1];
  assign _1736_ = _1735_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5765" *) _2265_;
  assign pout_mem_data_sel_1_last[1] = _1736_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5765" *) mem_re2_sel;
  assign _1737_ = _2682_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5766" *) mem_re_last_2d[2];
  assign _1738_ = _1737_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5766" *) _2265_;
  assign pout_mem_data_sel_1_last[2] = _1738_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5766" *) mem_re2_sel;
  assign _1739_ = _2682_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5767" *) mem_re_last_2d[3];
  assign _1740_ = _1739_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5767" *) _2265_;
  assign pout_mem_data_sel_1_last[3] = _1740_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5767" *) mem_re2_sel;
  assign _1741_ = _2682_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5768" *) mem_re_last_2d[4];
  assign _1742_ = _1741_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5768" *) _2266_;
  assign pout_mem_data_sel_1_last[4] = _1742_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5768" *) mem_re2_sel;
  assign _1743_ = _2682_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5769" *) mem_re_last_2d[5];
  assign _1744_ = _1743_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5769" *) _2266_;
  assign pout_mem_data_sel_1_last[5] = _1744_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5769" *) mem_re2_sel;
  assign _1745_ = _2682_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5770" *) mem_re_last_2d[6];
  assign _1746_ = _1745_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5770" *) _2266_;
  assign pout_mem_data_sel_1_last[6] = _1746_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5770" *) mem_re2_sel;
  assign _1747_ = _2682_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5771" *) mem_re_last_2d[7];
  assign _1748_ = _1747_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5771" *) _2266_;
  assign pout_mem_data_sel_1_last[7] = _1748_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5771" *) mem_re2_sel;
  assign pout_mem_data_sel_2_last[0] = _1734_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5773" *) mem_re3_sel;
  assign pout_mem_data_sel_2_last[1] = _1736_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5774" *) mem_re3_sel;
  assign _1749_ = _1737_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5775" *) _2266_;
  assign pout_mem_data_sel_2_last[2] = _1749_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5775" *) mem_re3_sel;
  assign _1750_ = _1739_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5776" *) _2266_;
  assign pout_mem_data_sel_2_last[3] = _1750_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5776" *) mem_re3_sel;
  assign _1751_ = _1741_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5777" *) _2267_;
  assign pout_mem_data_sel_2_last[4] = _1751_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5777" *) mem_re3_sel;
  assign _1752_ = _1743_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5778" *) _2267_;
  assign pout_mem_data_sel_2_last[5] = _1752_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5778" *) mem_re3_sel;
  assign _1753_ = _1745_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5779" *) _2268_;
  assign pout_mem_data_sel_2_last[6] = _1753_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5779" *) mem_re3_sel;
  assign _1754_ = _1747_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5780" *) _2268_;
  assign pout_mem_data_sel_2_last[7] = _1754_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5780" *) mem_re3_sel;
  assign pout_mem_data_sel_3_last[0] = _1734_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5782" *) mem_re4_sel;
  assign _1755_ = _1735_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5783" *) _2266_;
  assign pout_mem_data_sel_3_last[1] = _1755_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5783" *) mem_re4_sel;
  assign _1756_ = _1737_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5784" *) _2267_;
  assign pout_mem_data_sel_3_last[2] = _1756_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5784" *) mem_re4_sel;
  assign _1757_ = _1739_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5785" *) _2268_;
  assign pout_mem_data_sel_3_last[3] = _1757_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5785" *) mem_re4_sel;
  assign _1758_ = _1741_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5786" *) _2269_;
  assign pout_mem_data_sel_3_last[4] = _1758_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5786" *) mem_re4_sel;
  assign _1759_ = _1743_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5787" *) _2270_;
  assign pout_mem_data_sel_3_last[5] = _1759_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5787" *) mem_re4_sel;
  assign _1760_ = _1745_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5788" *) _2271_;
  assign pout_mem_data_sel_3_last[6] = _1760_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5788" *) mem_re4_sel;
  assign _1761_ = _1747_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5789" *) _2272_;
  assign pout_mem_data_sel_3_last[7] = _1761_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5789" *) mem_re4_sel;
  assign _1762_ = mem_data0_lst & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5791" *) { pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0], pout_mem_data_sel_last[0] };
  assign _1763_ = mem_data1_lst & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5792" *) { pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1], pout_mem_data_sel_last[1] };
  assign _1764_ = mem_data2_lst & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5793" *) { pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2], pout_mem_data_sel_last[2] };
  assign _1765_ = mem_data3_lst & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5794" *) { pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3], pout_mem_data_sel_last[3] };
  assign _1766_ = mem_data4_lst & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5795" *) { pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4], pout_mem_data_sel_last[4] };
  assign _1767_ = mem_data5_lst & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5796" *) { pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5], pout_mem_data_sel_last[5] };
  assign _1768_ = mem_data6_lst & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5797" *) { pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6], pout_mem_data_sel_last[6] };
  assign _1769_ = mem_data7_lst & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5798" *) { pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7], pout_mem_data_sel_last[7] };
  assign rd_line_out_done = wr_line_end_2d & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5805" *) rd_line_out;
  assign _1770_ = rd_line_out & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5816" *) _2273_;
  assign _1771_ = rd_sub_lbuf_end & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5828" *) _2274_;
  assign _1772_ = wr_surface_dat_done_2d & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5835" *) load_wr_stage2;
  assign _1773_ = rd_comb_lbuf_end & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5837" *) last_active_line_2d;
  assign _1774_ = _2275_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5841" *) rd_comb_lbuf_end;
  assign rd_lbuf_end = _1774_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5841" *) last_active_line_2d;
  assign _1775_ = load_wr_stage2 & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5845" *) _3113_;
  assign rd_pout_data_stage0 = load_wr_stage3_all & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5909" *) rd_pout_data_en_d;
  assign rd_pout_data_stage1_all = pout_data_stage1_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5983" *) pout_data_stage1_prdy;
  assign rd_pout_data_stage1 = rd_pout_data_stage1_all & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5984" *) rd_pout_data_en_2d;
  assign rd_pout_data_stage2_all = pout_data_stage2_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6057" *) pout_data_stage2_prdy;
  assign rd_pout_data_stage2 = rd_pout_data_stage2_all & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6058" *) rd_pout_data_en_3d;
  assign _1776_ = mem_re_2d & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6132" *) { load_wr_stage2, load_wr_stage2, load_wr_stage2, load_wr_stage2, load_wr_stage2, load_wr_stage2, load_wr_stage2, load_wr_stage2 };
  assign _1777_ = _1776_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6132" *) { mem_re1_sel, mem_re1_sel, mem_re1_sel, mem_re1_sel, mem_re1_sel, mem_re1_sel, mem_re1_sel, mem_re1_sel };
  assign pout_mem_data_sel_0 = _1777_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6132" *) { last_active_line_2d, last_active_line_2d, last_active_line_2d, last_active_line_2d, last_active_line_2d, last_active_line_2d, last_active_line_2d, last_active_line_2d };
  assign _1778_ = mem_re_2d[0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6134" *) load_wr_stage2;
  assign _1779_ = _1778_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6134" *) _2276_;
  assign _1780_ = _1779_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6134" *) last_active_line_2d;
  assign pout_mem_data_sel_1[0] = _1780_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6134" *) mem_re2_sel;
  assign _1781_ = mem_re_2d[1] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6135" *) load_wr_stage2;
  assign _1782_ = _1781_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6135" *) _2276_;
  assign _1783_ = _1782_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6135" *) last_active_line_2d;
  assign pout_mem_data_sel_1[1] = _1783_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6135" *) mem_re2_sel;
  assign _1784_ = mem_re_2d[2] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6136" *) load_wr_stage2;
  assign _1785_ = _1784_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6136" *) _2276_;
  assign _1786_ = _1785_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6136" *) last_active_line_2d;
  assign pout_mem_data_sel_1[2] = _1786_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6136" *) mem_re2_sel;
  assign _1787_ = mem_re_2d[3] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6137" *) load_wr_stage2;
  assign _1788_ = _1787_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6137" *) _2276_;
  assign _1789_ = _1788_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6137" *) last_active_line_2d;
  assign pout_mem_data_sel_1[3] = _1789_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6137" *) mem_re2_sel;
  assign _1790_ = mem_re_2d[4] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6138" *) load_wr_stage2;
  assign _1791_ = _1790_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6138" *) _2277_;
  assign _1792_ = _1791_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6138" *) last_active_line_2d;
  assign pout_mem_data_sel_1[4] = _1792_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6138" *) mem_re2_sel;
  assign _1793_ = mem_re_2d[5] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6139" *) load_wr_stage2;
  assign _1794_ = _1793_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6139" *) _2277_;
  assign _1795_ = _1794_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6139" *) last_active_line_2d;
  assign pout_mem_data_sel_1[5] = _1795_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6139" *) mem_re2_sel;
  assign _1796_ = mem_re_2d[6] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6140" *) load_wr_stage2;
  assign _1797_ = _1796_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6140" *) _2277_;
  assign _1798_ = _1797_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6140" *) last_active_line_2d;
  assign pout_mem_data_sel_1[6] = _1798_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6140" *) mem_re2_sel;
  assign _1799_ = mem_re_2d[7] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6141" *) load_wr_stage2;
  assign _1800_ = _1799_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6141" *) _2277_;
  assign _1801_ = _1800_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6141" *) last_active_line_2d;
  assign pout_mem_data_sel_1[7] = _1801_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6141" *) mem_re2_sel;
  assign pout_mem_data_sel_2[0] = _1780_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6143" *) mem_re3_sel;
  assign pout_mem_data_sel_2[1] = _1783_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6144" *) mem_re3_sel;
  assign _1802_ = _1784_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6145" *) _2277_;
  assign _1803_ = _1802_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6145" *) last_active_line_2d;
  assign pout_mem_data_sel_2[2] = _1803_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6145" *) mem_re3_sel;
  assign _1804_ = _1787_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6146" *) _2277_;
  assign _1805_ = _1804_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6146" *) last_active_line_2d;
  assign pout_mem_data_sel_2[3] = _1805_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6146" *) mem_re3_sel;
  assign _1806_ = _1790_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6147" *) _2278_;
  assign _1807_ = _1806_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6147" *) last_active_line_2d;
  assign pout_mem_data_sel_2[4] = _1807_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6147" *) mem_re3_sel;
  assign _1808_ = _1793_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6148" *) _2278_;
  assign _1809_ = _1808_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6148" *) last_active_line_2d;
  assign pout_mem_data_sel_2[5] = _1809_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6148" *) mem_re3_sel;
  assign _1810_ = _1796_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6149" *) _2279_;
  assign _1811_ = _1810_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6149" *) last_active_line_2d;
  assign pout_mem_data_sel_2[6] = _1811_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6149" *) mem_re3_sel;
  assign _1812_ = _1799_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6150" *) _2279_;
  assign _1813_ = _1812_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6150" *) last_active_line_2d;
  assign pout_mem_data_sel_2[7] = _1813_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6150" *) mem_re3_sel;
  assign pout_mem_data_sel_3[0] = _1780_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6152" *) mem_re4_sel;
  assign _1814_ = _1781_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6153" *) _2277_;
  assign _1815_ = _1814_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6153" *) last_active_line_2d;
  assign pout_mem_data_sel_3[1] = _1815_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6153" *) mem_re4_sel;
  assign _1816_ = _1784_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6154" *) _2278_;
  assign _1817_ = _1816_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6154" *) last_active_line_2d;
  assign pout_mem_data_sel_3[2] = _1817_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6154" *) mem_re4_sel;
  assign _1818_ = _1787_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6155" *) _2279_;
  assign _1819_ = _1818_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6155" *) last_active_line_2d;
  assign pout_mem_data_sel_3[3] = _1819_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6155" *) mem_re4_sel;
  assign _1820_ = _1790_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6156" *) _2280_;
  assign _1821_ = _1820_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6156" *) last_active_line_2d;
  assign pout_mem_data_sel_3[4] = _1821_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6156" *) mem_re4_sel;
  assign _1822_ = _1793_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6157" *) _2281_;
  assign _1823_ = _1822_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6157" *) last_active_line_2d;
  assign pout_mem_data_sel_3[5] = _1823_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6157" *) mem_re4_sel;
  assign _1824_ = _1796_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6158" *) _2282_;
  assign _1825_ = _1824_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6158" *) last_active_line_2d;
  assign pout_mem_data_sel_3[6] = _1825_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6158" *) mem_re4_sel;
  assign _1826_ = _1799_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6159" *) _2283_;
  assign _1827_ = _1826_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6159" *) last_active_line_2d;
  assign pout_mem_data_sel_3[7] = _1827_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6159" *) mem_re4_sel;
  assign padding_here = average_pooling_en & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6220" *) _2342_;
  assign _1828_ = _2435_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6325" *) average_pooling_en;
  assign _1829_ = data_hmult_16bit_0_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6374" *) _2436_;
  assign i16_less_neg_0_5_0 = data_hmult_16bit_0_ext[38] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6374" *) _2696_;
  assign _1830_ = data_hmult_16bit_1_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6375" *) _2438_;
  assign i16_less_neg_0_5_1 = data_hmult_16bit_1_ext[38] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6375" *) _2697_;
  assign _1831_ = data_hmult_16bit_2_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6376" *) _2440_;
  assign i16_less_neg_0_5_2 = data_hmult_16bit_2_ext[38] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6376" *) _2698_;
  assign _1832_ = data_hmult_16bit_3_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6377" *) _2442_;
  assign i16_less_neg_0_5_3 = data_hmult_16bit_3_ext[38] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6377" *) _2699_;
  assign _1833_ = data_hmult_16bit_0_ext[38] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6378" *) data_hmult_16bit_0_ext[15];
  assign i16_more_neg_0_5_0 = _1833_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6378" *) _3114_;
  assign _1834_ = data_hmult_16bit_1_ext[38] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6379" *) data_hmult_16bit_1_ext[15];
  assign i16_more_neg_0_5_1 = _1834_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6379" *) _3115_;
  assign _1835_ = data_hmult_16bit_2_ext[38] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6380" *) data_hmult_16bit_2_ext[15];
  assign i16_more_neg_0_5_2 = _1835_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6380" *) _3116_;
  assign _1836_ = data_hmult_16bit_3_ext[38] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6381" *) data_hmult_16bit_3_ext[15];
  assign i16_more_neg_0_5_3 = _1836_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6381" *) _3117_;
  assign _1837_ = data_hmult_8bit_0_lsb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6587" *) _2444_;
  assign i8_less_neg_0_5_0_l = data_hmult_8bit_0_lsb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6587" *) _2700_;
  assign _1838_ = data_hmult_8bit_0_msb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6588" *) _2446_;
  assign i8_less_neg_0_5_0_m = data_hmult_8bit_0_msb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6588" *) _2701_;
  assign _1839_ = data_hmult_8bit_1_lsb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6589" *) _2448_;
  assign i8_less_neg_0_5_1_l = data_hmult_8bit_1_lsb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6589" *) _2702_;
  assign _1840_ = data_hmult_8bit_1_msb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6590" *) _2450_;
  assign i8_less_neg_0_5_1_m = data_hmult_8bit_1_msb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6590" *) _2703_;
  assign _1841_ = data_hmult_8bit_2_lsb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6591" *) _2452_;
  assign i8_less_neg_0_5_2_l = data_hmult_8bit_2_lsb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6591" *) _2704_;
  assign _1842_ = data_hmult_8bit_2_msb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6592" *) _2454_;
  assign i8_less_neg_0_5_2_m = data_hmult_8bit_2_msb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6592" *) _2705_;
  assign _1843_ = data_hmult_8bit_3_lsb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6593" *) _2456_;
  assign i8_less_neg_0_5_3_l = data_hmult_8bit_3_lsb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6593" *) _2706_;
  assign _1844_ = data_hmult_8bit_3_msb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6594" *) _2458_;
  assign i8_less_neg_0_5_3_m = data_hmult_8bit_3_msb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6594" *) _2707_;
  assign _1845_ = data_hmult_8bit_0_lsb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6595" *) data_hmult_8bit_0_lsb_ext[15];
  assign i8_more_neg_0_5_0_l = _1845_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6595" *) _3118_;
  assign _1846_ = data_hmult_8bit_0_msb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6596" *) data_hmult_8bit_0_msb_ext[15];
  assign i8_more_neg_0_5_0_m = _1846_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6596" *) _3119_;
  assign _1847_ = data_hmult_8bit_1_lsb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6597" *) data_hmult_8bit_1_lsb_ext[15];
  assign i8_more_neg_0_5_1_l = _1847_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6597" *) _3120_;
  assign _1848_ = data_hmult_8bit_1_msb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6598" *) data_hmult_8bit_1_msb_ext[15];
  assign i8_more_neg_0_5_1_m = _1848_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6598" *) _3121_;
  assign _1849_ = data_hmult_8bit_2_lsb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6599" *) data_hmult_8bit_2_lsb_ext[15];
  assign i8_more_neg_0_5_2_l = _1849_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6599" *) _3122_;
  assign _1850_ = data_hmult_8bit_2_msb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6600" *) data_hmult_8bit_2_msb_ext[15];
  assign i8_more_neg_0_5_2_m = _1850_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6600" *) _3123_;
  assign _1851_ = data_hmult_8bit_3_lsb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6601" *) data_hmult_8bit_3_lsb_ext[15];
  assign i8_more_neg_0_5_3_l = _1851_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6601" *) _3124_;
  assign _1852_ = data_hmult_8bit_3_msb_ext[30] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6602" *) data_hmult_8bit_3_msb_ext[15];
  assign i8_more_neg_0_5_3_m = _1852_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6602" *) _3125_;
  assign _1853_ = data_vmult_16bit_0_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7029" *) _2460_;
  assign i16_vless_neg_0_5_0 = data_vmult_16bit_0_ext[35] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7029" *) _2708_;
  assign _1854_ = data_vmult_16bit_1_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7030" *) _2462_;
  assign i16_vless_neg_0_5_1 = data_vmult_16bit_1_ext[35] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7030" *) _2709_;
  assign _1855_ = data_vmult_16bit_2_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7031" *) _2464_;
  assign i16_vless_neg_0_5_2 = data_vmult_16bit_2_ext[35] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7031" *) _2710_;
  assign _1856_ = data_vmult_16bit_3_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7032" *) _2466_;
  assign i16_vless_neg_0_5_3 = data_vmult_16bit_3_ext[35] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7032" *) _2711_;
  assign _1857_ = data_vmult_16bit_0_ext[35] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7033" *) data_vmult_16bit_0_ext[15];
  assign i16_vmore_neg_0_5_0 = _1857_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7033" *) _3126_;
  assign _1858_ = data_vmult_16bit_1_ext[35] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7034" *) data_vmult_16bit_1_ext[15];
  assign i16_vmore_neg_0_5_1 = _1858_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7034" *) _3127_;
  assign _1859_ = data_vmult_16bit_2_ext[35] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7035" *) data_vmult_16bit_2_ext[15];
  assign i16_vmore_neg_0_5_2 = _1859_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7035" *) _3128_;
  assign _1860_ = data_vmult_16bit_3_ext[35] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7036" *) data_vmult_16bit_3_ext[15];
  assign i16_vmore_neg_0_5_3 = _1860_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7036" *) _3129_;
  assign _1861_ = data_vmult_8bit_0_lsb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7242" *) _2468_;
  assign i8_vless_neg_0_5_0_l = data_vmult_8bit_0_lsb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7242" *) _2712_;
  assign _1862_ = data_vmult_8bit_0_msb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7243" *) _2470_;
  assign i8_vless_neg_0_5_0_m = data_vmult_8bit_0_msb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7243" *) _2713_;
  assign _1863_ = data_vmult_8bit_1_lsb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7244" *) _2472_;
  assign i8_vless_neg_0_5_1_l = data_vmult_8bit_1_lsb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7244" *) _2714_;
  assign _1864_ = data_vmult_8bit_1_msb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7245" *) _2474_;
  assign i8_vless_neg_0_5_1_m = data_vmult_8bit_1_msb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7245" *) _2715_;
  assign _1865_ = data_vmult_8bit_2_lsb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7246" *) _2476_;
  assign i8_vless_neg_0_5_2_l = data_vmult_8bit_2_lsb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7246" *) _2716_;
  assign _1866_ = data_vmult_8bit_2_msb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7247" *) _2478_;
  assign i8_vless_neg_0_5_2_m = data_vmult_8bit_2_msb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7247" *) _2717_;
  assign _1867_ = data_vmult_8bit_3_lsb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7248" *) _2480_;
  assign i8_vless_neg_0_5_3_l = data_vmult_8bit_3_lsb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7248" *) _2718_;
  assign _1868_ = data_vmult_8bit_3_msb_ext[15] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7249" *) _2482_;
  assign i8_vless_neg_0_5_3_m = data_vmult_8bit_3_msb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7249" *) _2719_;
  assign _1869_ = data_vmult_8bit_0_lsb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7250" *) data_vmult_8bit_0_lsb_ext[15];
  assign i8_vmore_neg_0_5_0_l = _1869_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7250" *) _3130_;
  assign _1870_ = data_vmult_8bit_0_msb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7251" *) data_vmult_8bit_0_msb_ext[15];
  assign i8_vmore_neg_0_5_0_m = _1870_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7251" *) _3131_;
  assign _1871_ = data_vmult_8bit_1_lsb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7252" *) data_vmult_8bit_1_lsb_ext[15];
  assign i8_vmore_neg_0_5_1_l = _1871_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7252" *) _3132_;
  assign _1872_ = data_vmult_8bit_1_msb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7253" *) data_vmult_8bit_1_msb_ext[15];
  assign i8_vmore_neg_0_5_1_m = _1872_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7253" *) _3133_;
  assign _1873_ = data_vmult_8bit_2_lsb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7254" *) data_vmult_8bit_2_lsb_ext[15];
  assign i8_vmore_neg_0_5_2_l = _1873_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7254" *) _3134_;
  assign _1874_ = data_vmult_8bit_2_msb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7255" *) data_vmult_8bit_2_msb_ext[15];
  assign i8_vmore_neg_0_5_2_m = _1874_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7255" *) _3135_;
  assign _1875_ = data_vmult_8bit_3_lsb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7256" *) data_vmult_8bit_3_lsb_ext[15];
  assign i8_vmore_neg_0_5_3_l = _1875_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7256" *) _3136_;
  assign _1876_ = data_vmult_8bit_3_msb_ext[27] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7257" *) data_vmult_8bit_3_msb_ext[15];
  assign i8_vmore_neg_0_5_3_m = _1876_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7257" *) _3137_;
  assign int_dp2wdma_valid = pout_data_stage3_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7674" *) rd_pout_data_en_4d;
  assign fp16_add_in_rdy = din_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7781" *) _3016_;
  assign fp16_mean_pool_valid = fp16_mean_pool_cfg & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7783" *) wr_data_stage1_vld;
  assign _1877_ = fp16_mean_pool_valid & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7784" *) _3017_;
  assign fp16_4add_in_pvld[0] = _1877_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7784" *) din_rdy;
  assign _1878_ = fp16_mean_pool_valid & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7785" *) _3018_;
  assign fp16_4add_in_pvld[1] = _1878_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7785" *) din_rdy;
  assign _1879_ = fp16_mean_pool_valid & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7786" *) _3019_;
  assign fp16_4add_in_pvld[2] = _1879_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7786" *) din_rdy;
  assign _1880_ = fp16_mean_pool_valid & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7787" *) _3020_;
  assign fp16_4add_in_pvld[3] = _1880_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7787" *) din_rdy;
  assign _1881_ = fp16_mean_pool_valid & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7788" *) _3021_;
  assign fp16_4add_in_pvld[4] = _1881_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7788" *) din_rdy;
  assign _1882_ = fp16_mean_pool_valid & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7789" *) _3022_;
  assign fp16_4add_in_pvld[5] = _1882_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7789" *) din_rdy;
  assign _1883_ = fp16_mean_pool_valid & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7790" *) _3023_;
  assign fp16_4add_in_pvld[6] = _1883_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7790" *) din_rdy;
  assign _1884_ = fp16_mean_pool_valid & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7791" *) _3024_;
  assign fp16_4add_in_pvld[7] = _1884_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7791" *) din_rdy;
  assign din_vld_d0 = fp16_mean_pool_valid & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7792" *) _3016_;
  assign din_rdy_d4 = fp16_mul_pad_line_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7952" *) _3025_;
  assign _1885_ = fp16_mul_pad_line_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7953" *) _3026_;
  assign fp16_4add_out_prdy[0] = _1885_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7953" *) din_vld_d4;
  assign _1886_ = fp16_mul_pad_line_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7954" *) _3027_;
  assign fp16_4add_out_prdy[1] = _1886_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7954" *) din_vld_d4;
  assign _1887_ = fp16_mul_pad_line_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7955" *) _3028_;
  assign fp16_4add_out_prdy[2] = _1887_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7955" *) din_vld_d4;
  assign _1888_ = fp16_mul_pad_line_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7956" *) _3029_;
  assign fp16_4add_out_prdy[3] = _1888_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7956" *) din_vld_d4;
  assign _1889_ = fp16_mul_pad_line_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7957" *) _3030_;
  assign fp16_4add_out_prdy[4] = _1889_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7957" *) din_vld_d4;
  assign _1890_ = fp16_mul_pad_line_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7958" *) _3031_;
  assign fp16_4add_out_prdy[5] = _1890_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7958" *) din_vld_d4;
  assign _1891_ = fp16_mul_pad_line_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7959" *) _3032_;
  assign fp16_4add_out_prdy[6] = _1891_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7959" *) din_vld_d4;
  assign _1892_ = fp16_mul_pad_line_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7960" *) _3033_;
  assign fp16_4add_out_prdy[7] = _1892_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7960" *) din_vld_d4;
  assign fp_add_out_vld = din_vld_d4 & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7961" *) _3025_;
  assign _1893_ = fp_add_out_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7963" *) fp16_mul_pad_line_prdy;
  assign _1894_ = _1893_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7963" *) _2484_;
  assign fp_add_out_load = _1894_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7963" *) _2485_;
  assign fp_mem_we[0] = fp_add_out_load & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7968" *) din_pd_d4[246];
  assign fp_mem_we[1] = fp_add_out_load & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7973" *) din_pd_d4[247];
  assign fp_mem_we[2] = fp_add_out_load & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7978" *) din_pd_d4[248];
  assign fp_mem_we[3] = fp_add_out_load & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7983" *) din_pd_d4[249];
  assign fp_mem_we[4] = fp_add_out_load & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7988" *) din_pd_d4[250];
  assign fp_mem_we[5] = fp_add_out_load & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7993" *) din_pd_d4[251];
  assign fp_mem_we[6] = fp_add_out_load & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7998" *) din_pd_d4[252];
  assign fp_mem_we[7] = fp_add_out_load & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8003" *) din_pd_d4[253];
  assign _1895_ = { din_pd_d4[131:129], 11'b00000000000, fp_mem0_wdata[100:0] } & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8023" *) { din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121], din_pd_d4[121] };
  assign _1896_ = { din_pd_d4[135:133], 11'b00000000000, fp_mem1_wdata[100:0] } & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8024" *) { din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122], din_pd_d4[122] };
  assign _1897_ = { din_pd_d4[139:137], 11'b00000000000, fp_mem2_wdata[100:0] } & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8025" *) { din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123], din_pd_d4[123] };
  assign _1898_ = { din_pd_d4[143:141], 11'b00000000000, fp_mem3_wdata[100:0] } & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8026" *) { din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124], din_pd_d4[124] };
  assign _1899_ = { din_pd_d4[147:145], 11'b00000000000, fp_mem4_wdata[100:0] } & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8027" *) { din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125], din_pd_d4[125] };
  assign _1900_ = { din_pd_d4[151:149], 11'b00000000000, fp_mem5_wdata[100:0] } & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8028" *) { din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126], din_pd_d4[126] };
  assign _1901_ = { din_pd_d4[155:153], 11'b00000000000, fp_mem6_wdata[100:0] } & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8029" *) { din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127], din_pd_d4[127] };
  assign _1902_ = { din_pd_d4[159:157], 11'b00000000000, fp_mem7_wdata[100:0] } & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8030" *) { din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128], din_pd_d4[128] };
  assign _1903_ = din_pd_d4[114:0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8031" *) { din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161], din_pd_d4[161] };
  assign _1904_ = din_pd_d4[114:0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8032" *) { din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162], din_pd_d4[162] };
  assign _1905_ = din_pd_d4[114:0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8033" *) { din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163], din_pd_d4[163] };
  assign _1906_ = din_pd_d4[114:0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8034" *) { din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164], din_pd_d4[164] };
  assign _1907_ = din_pd_d4[114:0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8035" *) { din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165], din_pd_d4[165] };
  assign _1908_ = din_pd_d4[114:0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8036" *) { din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166], din_pd_d4[166] };
  assign _1909_ = din_pd_d4[114:0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8037" *) { din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167], din_pd_d4[167] };
  assign _1910_ = din_pd_d4[114:0] & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8038" *) { din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168], din_pd_d4[168] };
  assign fp16_mul_pad_line_prdy = _3034_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8787" *) fp16_mul_pad_line_in_rdy;
  assign _1911_ = fp16_mulw_in_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8788" *) fp16_mul_pad_line_rdy[1];
  assign fp16_mul_pad_line_vld[0] = _1911_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8788" *) fp16_mul_pad_line_in_rdy;
  assign _1912_ = fp16_mulw_in_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8789" *) fp16_mul_pad_line_rdy[0];
  assign fp16_mul_pad_line_vld[1] = _1912_ & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8789" *) fp16_mul_pad_line_in_rdy;
  assign fp16_mul_pad_line_in_vld_d0 = fp16_mulw_in_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8790" *) _3034_;
  assign fp16_mul_pad_line_in_rdy_d3 = fp_mulw_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8842" *) pad_line_sum_pvld;
  assign pad_line_sum_prdy = fp_mulw_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8843" *) fp16_mul_pad_line_in_vld_d3;
  assign fp16_mul_pad_line_pvld = pad_line_sum_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8844" *) fp16_mul_pad_line_in_vld_d3;
  assign fp16_add_pad_in_a_vld[0] = fp16_mul_pad_line_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8850" *) _3035_;
  assign fp16_add_pad_in_a_vld[1] = fp16_mul_pad_line_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8851" *) _3036_;
  assign fp16_add_pad_in_a_vld[2] = fp16_mul_pad_line_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8852" *) _3037_;
  assign fp16_add_pad_in_a_vld[3] = fp16_mul_pad_line_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8853" *) _3038_;
  assign fp16_add_pad_in_b_vld[0] = fp16_mul_pad_line_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8854" *) _3039_;
  assign fp16_add_pad_in_b_vld[1] = fp16_mul_pad_line_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8855" *) _3040_;
  assign fp16_add_pad_in_b_vld[2] = fp16_mul_pad_line_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8856" *) _3041_;
  assign fp16_add_pad_in_b_vld[3] = fp16_mul_pad_line_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8857" *) _3042_;
  assign fp16_add_pad_out_rdy[0] = fp16_mulw_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8910" *) _3043_;
  assign fp16_add_pad_out_rdy[1] = fp16_mulw_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8911" *) _3044_;
  assign fp16_add_pad_out_rdy[2] = fp16_mulw_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8912" *) _3045_;
  assign fp16_add_pad_out_rdy[3] = fp16_mulw_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8913" *) _3046_;
  assign fp16_mulw_in_a_vld[0] = fp16_add_pad_out_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8922" *) _3047_;
  assign fp16_mulw_in_a_vld[1] = fp16_add_pad_out_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8923" *) _3048_;
  assign fp16_mulw_in_a_vld[2] = fp16_add_pad_out_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8924" *) _3049_;
  assign fp16_mulw_in_a_vld[3] = fp16_add_pad_out_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8925" *) _3050_;
  assign fp16_mulw_in_b_vld[0] = fp16_add_pad_out_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8926" *) _3051_;
  assign fp16_mulw_in_b_vld[1] = fp16_add_pad_out_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8927" *) _3052_;
  assign fp16_mulw_in_b_vld[2] = fp16_add_pad_out_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8928" *) _3053_;
  assign fp16_mulw_in_b_vld[3] = fp16_add_pad_out_pvld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8929" *) _3054_;
  assign fp16_mulw_out_rdy[0] = fp16_mulv_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8983" *) _3055_;
  assign fp16_mulw_out_rdy[1] = fp16_mulv_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8984" *) _3056_;
  assign fp16_mulw_out_rdy[2] = fp16_mulv_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8985" *) _3057_;
  assign fp16_mulw_out_rdy[3] = fp16_mulv_rdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8986" *) _3058_;
  assign fp16_mulv_in_a_vld[0] = fp16_mulv_in_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8994" *) _3059_;
  assign fp16_mulv_in_a_vld[1] = fp16_mulv_in_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8995" *) _3060_;
  assign fp16_mulv_in_a_vld[2] = fp16_mulv_in_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8996" *) _3061_;
  assign fp16_mulv_in_a_vld[3] = fp16_mulv_in_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8997" *) _3062_;
  assign fp16_mulv_in_b_vld[0] = fp16_mulv_in_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8998" *) _3063_;
  assign fp16_mulv_in_b_vld[1] = fp16_mulv_in_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8999" *) _3064_;
  assign fp16_mulv_in_b_vld[2] = fp16_mulv_in_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9000" *) _3065_;
  assign fp16_mulv_in_b_vld[3] = fp16_mulv_in_vld & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9001" *) _3066_;
  assign fp17T16_out_rdy[0] = fp_dp2wdma_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9099" *) _3067_;
  assign fp17T16_out_rdy[1] = fp_dp2wdma_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9100" *) _3068_;
  assign fp17T16_out_rdy[2] = fp_dp2wdma_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9101" *) _3069_;
  assign fp17T16_out_rdy[3] = fp_dp2wdma_prdy & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9102" *) _3070_;
  assign fp_dp2wdma_prdy = fp16_mean_pool_cfg & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9105" *) pdp_dp2wdma_ready;
  assign average_pooling_en = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1144" *) pooling_type_cfg;
  assign int8_en = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1145" *) reg2dp_input_data;
  assign data_c_end = c_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1156" *) 2'b11;
  assign _2011_ = wr_line_dat_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1168" *) pout_width_cur;
  assign last_line_in = wr_surface_dat_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1180" *) reg2dp_cube_in_height;
  assign _2012_ = { _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[9:0] } == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1201" *) surface_cnt_rd;
  assign _2013_ = wr_splitc_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1213" *) pooling_splitw_num_cfg;
  assign _2014_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1218" *) wr_splitc_cnt;
  assign _2015_ = strip_ycnt_stride == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1302" *) pooling_stride_v_cfg;
  assign _2017_ = pad_r_remain == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1465" *) stride_6x;
  assign _2018_ = pad_r_remain == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1467" *) stride_5x;
  assign _2019_ = pad_r_remain == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1469" *) { pooling_stride_v, 2'b00 };
  assign _2020_ = pad_r_remain == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1471" *) stride_3x;
  assign _2021_ = pad_r_remain == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1473" *) { pooling_stride_v, 1'b0 };
  assign _1228_ = pad_r_remain == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1475" *) pooling_stride_v;
  assign _2022_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1486" *) flush_num_cal;
  assign _2023_ = flush_in_next_surf == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1562" *) 2'b10;
  assign _2024_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1563" *) bubble_num;
  assign _2025_ = bubble_num == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1566" *) 1'b1;
  assign _2026_ = bubble_num == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1569" *) 2'b10;
  assign _2027_ = bubble_num == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1572" *) 2'b11;
  assign _2028_ = bubble_num == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1575" *) 3'b100;
  assign _2029_ = flush_in_next_surf == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1598" *) 2'b11;
  assign _2030_ = flush_in_next_surf == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1637" *) 3'b100;
  assign _2031_ = flush_in_next_surf == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1677" *) 3'b101;
  assign _2032_ = flush_in_next_surf == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1716" *) 3'b110;
  assign _2033_ = flush_in_next_surf == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1751" *) 3'b111;
  assign _2034_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) next2_1;
  assign _2035_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) next2_1;
  assign _2036_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) next2_1;
  assign _2037_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) next2_1;
  assign _2038_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) next2_1;
  assign _2039_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) next2_1;
  assign _2040_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *) next2_0;
  assign _2041_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *) next2_0;
  assign _2042_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *) next2_0;
  assign _2043_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *) next2_0;
  assign _2044_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *) next2_0;
  assign _2045_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *) next2_0;
  assign _2046_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) next3_2;
  assign _2047_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) next3_2;
  assign _2048_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) next3_2;
  assign _2049_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) next3_2;
  assign _2050_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) next3_2;
  assign _2051_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) next3_2;
  assign _2052_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) next3_1;
  assign _2053_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) next3_1;
  assign _2054_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) next3_1;
  assign _2055_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) next3_1;
  assign _2056_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) next3_1;
  assign _2057_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) next3_1;
  assign _2058_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *) next3_0;
  assign _2059_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *) next3_0;
  assign _2060_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *) next3_0;
  assign _2061_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *) next3_0;
  assign _2062_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *) next3_0;
  assign _2063_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *) next3_0;
  assign _2064_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) next4_3;
  assign _2065_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) next4_3;
  assign _2066_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) next4_3;
  assign _2067_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) next4_3;
  assign _2068_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) next4_3;
  assign _2069_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) next4_3;
  assign _2070_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) next4_2;
  assign _2071_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) next4_2;
  assign _2072_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) next4_2;
  assign _2073_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) next4_2;
  assign _2074_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) next4_2;
  assign _2075_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) next4_2;
  assign _2076_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) next4_1;
  assign _2077_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) next4_1;
  assign _2078_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) next4_1;
  assign _2079_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) next4_1;
  assign _2080_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) next4_1;
  assign _2081_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) next4_1;
  assign _2082_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *) next4_0;
  assign _2083_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *) next4_0;
  assign _2084_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *) next4_0;
  assign _2085_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *) next4_0;
  assign _2086_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *) next4_0;
  assign _2087_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *) next4_0;
  assign _2088_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) next5_4;
  assign _2089_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) next5_4;
  assign _2090_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) next5_4;
  assign _2091_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) next5_4;
  assign _2092_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) next5_4;
  assign _2093_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) next5_4;
  assign _2094_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) next5_3;
  assign _2095_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) next5_3;
  assign _2096_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) next5_3;
  assign _2097_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) next5_3;
  assign _2098_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) next5_3;
  assign _2099_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) next5_3;
  assign _2100_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) next5_2;
  assign _2101_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) next5_2;
  assign _2102_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) next5_2;
  assign _2103_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) next5_2;
  assign _2104_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) next5_2;
  assign _2105_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) next5_2;
  assign _2106_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) next5_1;
  assign _2107_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) next5_1;
  assign _2108_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) next5_1;
  assign _2109_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) next5_1;
  assign _2110_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) next5_1;
  assign _2111_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) next5_1;
  assign _2112_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *) next5_0;
  assign _2113_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *) next5_0;
  assign _2114_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *) next5_0;
  assign _2115_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *) next5_0;
  assign _2116_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *) next5_0;
  assign _2117_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *) next5_0;
  assign _2118_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) next6_5;
  assign _2119_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) next6_5;
  assign _2120_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) next6_5;
  assign _2121_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) next6_5;
  assign _2122_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) next6_5;
  assign _2123_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) next6_5;
  assign _2124_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) next6_4;
  assign _2125_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) next6_4;
  assign _2126_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) next6_4;
  assign _2127_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) next6_4;
  assign _2128_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) next6_4;
  assign _2129_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) next6_4;
  assign _2130_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) next6_3;
  assign _2131_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) next6_3;
  assign _2132_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) next6_3;
  assign _2133_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) next6_3;
  assign _2134_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) next6_3;
  assign _2135_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) next6_3;
  assign _2136_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) next6_2;
  assign _2137_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) next6_2;
  assign _2138_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) next6_2;
  assign _2139_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) next6_2;
  assign _2140_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) next6_2;
  assign _2141_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) next6_2;
  assign _2142_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) next6_1;
  assign _2143_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) next6_1;
  assign _2144_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) next6_1;
  assign _2145_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) next6_1;
  assign _2146_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) next6_1;
  assign _2147_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) next6_1;
  assign _2148_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *) next6_0;
  assign _2149_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *) next6_0;
  assign _2150_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *) next6_0;
  assign _2151_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *) next6_0;
  assign _2152_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *) next6_0;
  assign _2153_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *) next6_0;
  assign _2154_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) next7_6;
  assign _2155_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) next7_6;
  assign _2156_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) next7_6;
  assign _2157_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) next7_6;
  assign _2158_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) next7_6;
  assign _2159_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) next7_6;
  assign _2160_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) next7_5;
  assign _2161_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) next7_5;
  assign _2162_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) next7_5;
  assign _2163_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) next7_5;
  assign _2164_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) next7_5;
  assign _2165_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) next7_5;
  assign _2166_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) next7_4;
  assign _2167_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) next7_4;
  assign _2168_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) next7_4;
  assign _2169_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) next7_4;
  assign _2170_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) next7_4;
  assign _2171_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) next7_4;
  assign _2172_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) next7_3;
  assign _2173_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) next7_3;
  assign _2174_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) next7_3;
  assign _2175_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) next7_3;
  assign _2176_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) next7_3;
  assign _2177_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) next7_3;
  assign _2178_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) next7_2;
  assign _2179_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) next7_2;
  assign _2180_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) next7_2;
  assign _2181_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) next7_2;
  assign _2182_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) next7_2;
  assign _2183_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) next7_2;
  assign _2184_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) next7_1;
  assign _2185_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) next7_1;
  assign _2186_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) next7_1;
  assign _2187_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) next7_1;
  assign _2188_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) next7_1;
  assign _2189_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) next7_1;
  assign _2190_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *) next7_0;
  assign _2191_ = up_pnum1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *) next7_0;
  assign _2192_ = up_pnum2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *) next7_0;
  assign _2193_ = up_pnum3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *) next7_0;
  assign _2194_ = up_pnum4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *) next7_0;
  assign _2195_ = up_pnum5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *) next7_0;
  assign unit2d_cnt_pooling_end = unit2d_cnt_pooling == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1862" *) unit2d_cnt_pooling_max;
  assign _2196_ = unit2d_cnt_pooling_a1 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1870" *) unit2d_cnt_pooling_max;
  assign _2197_ = unit2d_cnt_pooling_a2 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1878" *) unit2d_cnt_pooling_max;
  assign _2198_ = unit2d_cnt_pooling_a3 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1886" *) unit2d_cnt_pooling_max;
  assign _2199_ = unit2d_cnt_pooling_a4 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1894" *) unit2d_cnt_pooling_max;
  assign _2200_ = unit2d_cnt_pooling_a5 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1902" *) unit2d_cnt_pooling_max;
  assign _2201_ = unit2d_cnt_pooling_a6 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1910" *) unit2d_cnt_pooling_max;
  assign _2202_ = unit2d_cnt_pooling_a7 == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1918" *) unit2d_cnt_pooling_max;
  assign _2203_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1934" *) padding_v_cfg;
  assign _2204_ = padding_v_cfg == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1940" *) 1'b1;
  assign _2205_ = pooling_stride_v == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1941" *) 1'b1;
  assign _2206_ = padding_v_cfg == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1954" *) 2'b10;
  assign _2207_ = pooling_stride_v == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1961" *) 2'b10;
  assign _2208_ = padding_v_cfg == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1974" *) 2'b11;
  assign _2209_ = pooling_stride_v == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1981" *) 2'b11;
  assign _2210_ = padding_v_cfg == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1994" *) 3'b100;
  assign _2211_ = pooling_stride_v == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2007" *) 3'b100;
  assign _2212_ = padding_v_cfg == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2020" *) 3'b101;
  assign _2213_ = pooling_stride_v == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2033" *) 3'b101;
  assign _2214_ = channel_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2117" *) 2'b11;
  assign _2215_ = line_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2131" *) pout_width_cur_latch;
  assign _2216_ = bubble_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2145" *) bubble_num_dec;
  assign _2217_ = last_out_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2182" *) first_out_num_dec2;
  assign _2218_ = last_out_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2182" *) flush_num_dec1;
  assign _2219_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2252" *) reg2dp_cube_out_width;
  assign _2220_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2254" *) reg2dp_partial_width_out_first;
  assign _2221_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2256" *) reg2dp_partial_width_out_last;
  assign _2222_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2258" *) reg2dp_partial_width_out_mid;
  assign _2223_ = one_width_bubble_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2285" *) 2'b10;
  assign _2224_ = strip_ycnt_psize == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2287" *) pooling_size_v_cfg;
  assign stride_trig_end = unit2d_cnt_pooling_max == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2306" *) unit2d_cnt_stride;
  assign _2225_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2334" *) unit2d_cnt_pooling;
  assign _2226_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2348" *) unit2d_cnt_stride;
  assign _2227_ = unit2d_cnt_pooling == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2350" *) 1'b1;
  assign _2228_ = unit2d_cnt_stride == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2364" *) 1'b1;
  assign _2229_ = unit2d_cnt_pooling == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2366" *) 2'b10;
  assign _2230_ = unit2d_cnt_stride == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2380" *) 2'b10;
  assign _2231_ = unit2d_cnt_pooling == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2382" *) 2'b11;
  assign _2232_ = unit2d_cnt_stride == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2396" *) 2'b11;
  assign _2233_ = unit2d_cnt_pooling == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2398" *) 3'b100;
  assign _2234_ = unit2d_cnt_stride == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2412" *) 3'b100;
  assign _2235_ = unit2d_cnt_pooling == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2414" *) 3'b101;
  assign _2236_ = unit2d_cnt_stride == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2428" *) 3'b101;
  assign _2237_ = unit2d_cnt_pooling == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2430" *) 3'b110;
  assign _2238_ = unit2d_cnt_stride == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2444" *) 3'b110;
  assign _2239_ = unit2d_cnt_pooling == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2446" *) 3'b111;
  assign _2240_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3327" *) wr_sub_lbuf_cnt;
  assign _2241_ = wr_sub_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3328" *) 1'b1;
  assign _2242_ = wr_sub_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3329" *) 2'b10;
  assign _2243_ = wr_sub_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3330" *) 2'b11;
  assign _2244_ = wr_sub_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3331" *) 3'b100;
  assign _2245_ = wr_sub_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3332" *) 3'b101;
  assign _2246_ = wr_sub_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3333" *) 3'b110;
  assign _2247_ = wr_sub_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3334" *) 3'b111;
  assign _1051_ = buffer_lines_num == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3403" *) 1'b1;
  assign _1052_ = buffer_lines_num == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3404" *) 2'b10;
  assign _2248_ = buffer_lines_num == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3405" *) 2'b11;
  assign _2249_ = buffer_lines_num == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3405" *) 3'b100;
  assign _2250_ = { _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[3:0] } == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3426" *) wr_sub_lbuf_cnt;
  assign _2251_ = sub_lbuf_dout_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3440" *) 6'b111111;
  assign _0980_ = pooling_type_cfg == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3583" *) 2'b10;
  assign _0979_ = pooling_type_cfg == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3584" *) 1'b1;
  assign unit2d_cnt_pooling_last_end = unit2d_cnt_pooling_last == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5049" *) unit2d_cnt_pooling_max;
  assign _2253_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5053" *) unit2d_cnt_pooling_last;
  assign _2254_ = unit2d_cnt_pooling_last == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5054" *) 1'b1;
  assign _2255_ = unit2d_cnt_pooling_last == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5055" *) 2'b10;
  assign _2256_ = unit2d_cnt_pooling_last == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5056" *) 2'b11;
  assign _2257_ = unit2d_cnt_pooling_last == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5057" *) 3'b100;
  assign _2258_ = unit2d_cnt_pooling_last == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5058" *) 3'b101;
  assign _2259_ = unit2d_cnt_pooling_last == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5059" *) 3'b110;
  assign _2260_ = unit2d_cnt_pooling_last == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5060" *) 3'b111;
  assign _2265_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5764" *) unit2d_cnt_pooling_last_2d;
  assign _2266_ = unit2d_cnt_pooling_last_2d == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5768" *) 1'b1;
  assign _2267_ = unit2d_cnt_pooling_last_2d == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5777" *) 2'b10;
  assign _2268_ = unit2d_cnt_pooling_last_2d == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5779" *) 2'b11;
  assign _2269_ = unit2d_cnt_pooling_last_2d == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5786" *) 3'b100;
  assign _2270_ = unit2d_cnt_pooling_last_2d == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5787" *) 3'b101;
  assign _2271_ = unit2d_cnt_pooling_last_2d == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5788" *) 3'b110;
  assign _2272_ = unit2d_cnt_pooling_last_2d == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5789" *) 3'b111;
  assign _2273_ = rd_line_out_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5816" *) 6'b111111;
  assign _2274_ = rd_sub_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5828" *) { _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[3:0] };
  assign _2275_ = rd_comb_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5841" *) { _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[3:0] };
  assign _2276_ = ! (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6134" *) rd_comb_lbuf_cnt;
  assign _2277_ = rd_comb_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6138" *) 1'b1;
  assign _2278_ = rd_comb_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6147" *) 2'b10;
  assign _2279_ = rd_comb_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6149" *) 2'b11;
  assign _2280_ = rd_comb_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6156" *) 3'b100;
  assign _2281_ = rd_comb_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6157" *) 3'b101;
  assign _2282_ = rd_comb_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6158" *) 3'b110;
  assign _2283_ = rd_comb_lbuf_cnt == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6159" *) 3'b111;
  assign fp16_en = reg2dp_input_data == (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8921" *) 2'b10;
  assign _2284_ = 3'b101 >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1236" *) pooling_size_v_cfg;
  assign pooling_stride_big = pooling_stride_v_cfg >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1239" *) pooling_size_v_cfg;
  assign _2285_ = padding_v_cfg >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1279" *) 3'b110;
  assign _2286_ = padding_v_cfg >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1280" *) 2'b11;
  assign _2287_ = pooling_size_v_cfg >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1390" *) pooling_stride_v_cfg;
  assign _2288_ = flush_num >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1520" *) first_out_num;
  assign _2289_ = padding_stride_num >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2331" *) 1'b0;
  assign _2290_ = padding_stride_num >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2347" *) 1'b1;
  assign _2291_ = padding_stride_num >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2363" *) 2'b10;
  assign _2292_ = padding_stride_num >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2379" *) 2'b11;
  assign _2293_ = padding_stride_num >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2395" *) 3'b100;
  assign _2294_ = padding_stride_num >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2411" *) 3'b101;
  assign _2295_ = padding_stride_num >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2427" *) 3'b110;
  assign _2296_ = padding_stride_num >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2443" *) 3'b111;
  assign _1056_ = buffer_lines_num >= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3406" *) 3'b101;
  assign padding_stride4_num[0] = padding_v_cfg > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1282" *) pooling_stride_v_cfg;
  assign _2297_ = pooling_splitw_num_cfg > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2258" *) 1'b1;
  assign _0403_ = $signed(_0002_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0000_);
  assign _0467_ = $signed(_0102_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0100_);
  assign _0531_ = $signed(_0202_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0200_);
  assign _0595_ = $signed(_0302_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0300_);
  assign _0411_ = $signed(_0016_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0000_);
  assign _0475_ = $signed(_0116_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0100_);
  assign _0539_ = $signed(_0216_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0200_);
  assign _0603_ = $signed(_0316_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0300_);
  assign _0419_ = $signed(_0028_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0000_);
  assign _0483_ = $signed(_0128_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0100_);
  assign _0547_ = $signed(_0228_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0200_);
  assign _0611_ = $signed(_0328_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0300_);
  assign _0427_ = $signed(_0040_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0000_);
  assign _0491_ = $signed(_0140_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0100_);
  assign _0555_ = $signed(_0240_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0200_);
  assign _0619_ = $signed(_0340_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0300_);
  assign _0435_ = $signed(_0052_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0000_);
  assign _0499_ = $signed(_0152_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0100_);
  assign _0563_ = $signed(_0252_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0200_);
  assign _0627_ = $signed(_0352_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0300_);
  assign _0443_ = $signed(_0064_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0000_);
  assign _0507_ = $signed(_0164_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0100_);
  assign _0571_ = $signed(_0264_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0200_);
  assign _0635_ = $signed(_0364_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0300_);
  assign _0451_ = $signed(_0076_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0000_);
  assign _0515_ = $signed(_0176_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0100_);
  assign _0579_ = $signed(_0276_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0200_);
  assign _0643_ = $signed(_0376_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0300_);
  assign _0459_ = $signed(_0088_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0000_);
  assign _0523_ = $signed(_0188_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0100_);
  assign _0587_ = $signed(_0288_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0200_);
  assign _0651_ = $signed(_0388_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3478" *) $signed(_0300_);
  assign _0405_ = $signed(_0003_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0001_);
  assign _0469_ = $signed(_0103_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0101_);
  assign _0533_ = $signed(_0203_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0201_);
  assign _0597_ = $signed(_0303_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0301_);
  assign _0413_ = $signed(_0017_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0001_);
  assign _0477_ = $signed(_0117_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0101_);
  assign _0541_ = $signed(_0217_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0201_);
  assign _0605_ = $signed(_0317_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0301_);
  assign _0421_ = $signed(_0029_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0001_);
  assign _0485_ = $signed(_0129_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0101_);
  assign _0549_ = $signed(_0229_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0201_);
  assign _0613_ = $signed(_0329_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0301_);
  assign _0429_ = $signed(_0041_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0001_);
  assign _0493_ = $signed(_0141_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0101_);
  assign _0557_ = $signed(_0241_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0201_);
  assign _0621_ = $signed(_0341_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0301_);
  assign _0437_ = $signed(_0053_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0001_);
  assign _0501_ = $signed(_0153_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0101_);
  assign _0565_ = $signed(_0253_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0201_);
  assign _0629_ = $signed(_0353_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0301_);
  assign _0445_ = $signed(_0065_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0001_);
  assign _0509_ = $signed(_0165_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0101_);
  assign _0573_ = $signed(_0265_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0201_);
  assign _0637_ = $signed(_0365_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0301_);
  assign _0453_ = $signed(_0077_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0001_);
  assign _0517_ = $signed(_0177_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0101_);
  assign _0581_ = $signed(_0277_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0201_);
  assign _0645_ = $signed(_0377_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0301_);
  assign _0461_ = $signed(_0089_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0001_);
  assign _0525_ = $signed(_0189_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0101_);
  assign _0589_ = $signed(_0289_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0201_);
  assign _0653_ = $signed(_0389_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3479" *) $signed(_0301_);
  assign _0401_ = $signed(_0007_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0006_);
  assign _0465_ = $signed(_0107_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0106_);
  assign _0529_ = $signed(_0207_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0206_);
  assign _0593_ = $signed(_0307_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0306_);
  assign _0409_ = $signed(_0019_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0006_);
  assign _0473_ = $signed(_0119_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0106_);
  assign _0537_ = $signed(_0219_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0206_);
  assign _0601_ = $signed(_0319_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0306_);
  assign _0417_ = $signed(_0031_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0006_);
  assign _0481_ = $signed(_0131_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0106_);
  assign _0545_ = $signed(_0231_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0206_);
  assign _0609_ = $signed(_0331_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0306_);
  assign _0425_ = $signed(_0043_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0006_);
  assign _0489_ = $signed(_0143_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0106_);
  assign _0553_ = $signed(_0243_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0206_);
  assign _0617_ = $signed(_0343_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0306_);
  assign _0433_ = $signed(_0055_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0006_);
  assign _0497_ = $signed(_0155_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0106_);
  assign _0561_ = $signed(_0255_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0206_);
  assign _0625_ = $signed(_0355_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0306_);
  assign _0441_ = $signed(_0067_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0006_);
  assign _0505_ = $signed(_0167_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0106_);
  assign _0569_ = $signed(_0267_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0206_);
  assign _0633_ = $signed(_0367_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0306_);
  assign _0449_ = $signed(_0079_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0006_);
  assign _0513_ = $signed(_0179_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0106_);
  assign _0577_ = $signed(_0279_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0206_);
  assign _0641_ = $signed(_0379_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0306_);
  assign _0457_ = $signed(_0091_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0006_);
  assign _0521_ = $signed(_0191_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0106_);
  assign _0585_ = $signed(_0291_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0206_);
  assign _0649_ = $signed(_0391_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3480" *) $signed(_0306_);
  assign _2298_ = _0004_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0005_[14:0];
  assign _2299_ = _0104_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0105_[14:0];
  assign _2300_ = _0204_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0205_[14:0];
  assign _2301_ = _0304_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0305_[14:0];
  assign _2302_ = _0004_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0018_[14:0];
  assign _2303_ = _0104_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0118_[14:0];
  assign _2304_ = _0204_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0218_[14:0];
  assign _2305_ = _0304_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0318_[14:0];
  assign _2306_ = _0004_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0030_[14:0];
  assign _2307_ = _0104_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0130_[14:0];
  assign _2308_ = _0204_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0230_[14:0];
  assign _2309_ = _0304_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0330_[14:0];
  assign _2310_ = _0004_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0042_[14:0];
  assign _2311_ = _0104_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0142_[14:0];
  assign _2312_ = _0204_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0242_[14:0];
  assign _2313_ = _0304_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0342_[14:0];
  assign _2314_ = _0004_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0054_[14:0];
  assign _2315_ = _0104_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0154_[14:0];
  assign _2316_ = _0204_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0254_[14:0];
  assign _2317_ = _0304_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0354_[14:0];
  assign _2318_ = _0004_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0066_[14:0];
  assign _2319_ = _0104_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0166_[14:0];
  assign _2320_ = _0204_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0266_[14:0];
  assign _2321_ = _0304_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0366_[14:0];
  assign _2322_ = _0004_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0078_[14:0];
  assign _2323_ = _0104_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0178_[14:0];
  assign _2324_ = _0204_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0278_[14:0];
  assign _2325_ = _0304_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0378_[14:0];
  assign _2326_ = _0004_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0090_[14:0];
  assign _2327_ = _0104_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0190_[14:0];
  assign _2328_ = _0204_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0290_[14:0];
  assign _2329_ = _0304_[14:0] > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0390_[14:0];
  assign _0011_ = $signed(_0000_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0002_);
  assign _0111_ = $signed(_0100_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0102_);
  assign _0211_ = $signed(_0200_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0202_);
  assign _0311_ = $signed(_0300_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0302_);
  assign _0023_ = $signed(_0000_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0016_);
  assign _0123_ = $signed(_0100_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0116_);
  assign _0223_ = $signed(_0200_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0216_);
  assign _0323_ = $signed(_0300_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0316_);
  assign _0035_ = $signed(_0000_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0028_);
  assign _0135_ = $signed(_0100_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0128_);
  assign _0235_ = $signed(_0200_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0228_);
  assign _0335_ = $signed(_0300_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0328_);
  assign _0047_ = $signed(_0000_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0040_);
  assign _0147_ = $signed(_0100_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0140_);
  assign _0247_ = $signed(_0200_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0240_);
  assign _0347_ = $signed(_0300_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0340_);
  assign _0059_ = $signed(_0000_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0052_);
  assign _0159_ = $signed(_0100_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0152_);
  assign _0259_ = $signed(_0200_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0252_);
  assign _0359_ = $signed(_0300_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0352_);
  assign _0071_ = $signed(_0000_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0064_);
  assign _0171_ = $signed(_0100_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0164_);
  assign _0271_ = $signed(_0200_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0264_);
  assign _0371_ = $signed(_0300_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0364_);
  assign _0083_ = $signed(_0000_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0076_);
  assign _0183_ = $signed(_0100_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0176_);
  assign _0283_ = $signed(_0200_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0276_);
  assign _0383_ = $signed(_0300_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0376_);
  assign _0095_ = $signed(_0000_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0088_);
  assign _0195_ = $signed(_0100_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0188_);
  assign _0295_ = $signed(_0200_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0288_);
  assign _0395_ = $signed(_0300_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3520" *) $signed(_0388_);
  assign _0013_ = $signed(_0001_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0003_);
  assign _0113_ = $signed(_0101_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0103_);
  assign _0213_ = $signed(_0201_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0203_);
  assign _0313_ = $signed(_0301_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0303_);
  assign _0025_ = $signed(_0001_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0017_);
  assign _0125_ = $signed(_0101_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0117_);
  assign _0225_ = $signed(_0201_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0217_);
  assign _0325_ = $signed(_0301_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0317_);
  assign _0037_ = $signed(_0001_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0029_);
  assign _0137_ = $signed(_0101_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0129_);
  assign _0237_ = $signed(_0201_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0229_);
  assign _0337_ = $signed(_0301_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0329_);
  assign _0049_ = $signed(_0001_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0041_);
  assign _0149_ = $signed(_0101_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0141_);
  assign _0249_ = $signed(_0201_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0241_);
  assign _0349_ = $signed(_0301_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0341_);
  assign _0061_ = $signed(_0001_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0053_);
  assign _0161_ = $signed(_0101_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0153_);
  assign _0261_ = $signed(_0201_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0253_);
  assign _0361_ = $signed(_0301_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0353_);
  assign _0073_ = $signed(_0001_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0065_);
  assign _0173_ = $signed(_0101_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0165_);
  assign _0273_ = $signed(_0201_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0265_);
  assign _0373_ = $signed(_0301_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0365_);
  assign _0085_ = $signed(_0001_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0077_);
  assign _0185_ = $signed(_0101_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0177_);
  assign _0285_ = $signed(_0201_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0277_);
  assign _0385_ = $signed(_0301_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0377_);
  assign _0097_ = $signed(_0001_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0089_);
  assign _0197_ = $signed(_0101_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0189_);
  assign _0297_ = $signed(_0201_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0289_);
  assign _0397_ = $signed(_0301_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3521" *) $signed(_0389_);
  assign _0009_ = $signed(_0006_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0007_);
  assign _0109_ = $signed(_0106_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0107_);
  assign _0209_ = $signed(_0206_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0207_);
  assign _0309_ = $signed(_0306_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0307_);
  assign _0021_ = $signed(_0006_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0019_);
  assign _0121_ = $signed(_0106_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0119_);
  assign _0221_ = $signed(_0206_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0219_);
  assign _0321_ = $signed(_0306_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0319_);
  assign _0033_ = $signed(_0006_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0031_);
  assign _0133_ = $signed(_0106_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0131_);
  assign _0233_ = $signed(_0206_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0231_);
  assign _0333_ = $signed(_0306_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0331_);
  assign _0045_ = $signed(_0006_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0043_);
  assign _0145_ = $signed(_0106_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0143_);
  assign _0245_ = $signed(_0206_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0243_);
  assign _0345_ = $signed(_0306_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0343_);
  assign _0057_ = $signed(_0006_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0055_);
  assign _0157_ = $signed(_0106_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0155_);
  assign _0257_ = $signed(_0206_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0255_);
  assign _0357_ = $signed(_0306_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0355_);
  assign _0069_ = $signed(_0006_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0067_);
  assign _0169_ = $signed(_0106_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0167_);
  assign _0269_ = $signed(_0206_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0267_);
  assign _0369_ = $signed(_0306_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0367_);
  assign _0081_ = $signed(_0006_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0079_);
  assign _0181_ = $signed(_0106_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0179_);
  assign _0281_ = $signed(_0206_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0279_);
  assign _0381_ = $signed(_0306_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0379_);
  assign _0093_ = $signed(_0006_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0091_);
  assign _0193_ = $signed(_0106_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0191_);
  assign _0293_ = $signed(_0206_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0291_);
  assign _0393_ = $signed(_0306_) > (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3522" *) $signed(_0391_);
  assign _2330_ = strip_ycnt_stride_f <= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1396" *) pooling_size_v_cfg;
  assign last_pooling_flag = rest_height_use <= (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2328" *) pooling_size_v_cfg;
  assign _2331_ = _1289_ || (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2098" *) _1291_;
  assign _2332_ = reg2dp_pad_bottom_cfg < (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1422" *) pooling_stride_v;
  assign _2333_ = reg2dp_pad_bottom_cfg < (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1424" *) { pooling_stride_v, 1'b0 };
  assign _2334_ = reg2dp_pad_bottom_cfg < (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1426" *) stride_3x;
  assign _2335_ = reg2dp_pad_bottom_cfg < (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1428" *) { pooling_stride_v, 2'b00 };
  assign _2336_ = reg2dp_pad_bottom_cfg < (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1430" *) stride_5x;
  assign _2337_ = reg2dp_pad_bottom_cfg < (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1432" *) stride_6x;
  assign _2338_ = reg2dp_pad_bottom_cfg < (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1434" *) stride_7x;
  assign _2339_ = h_pt < (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1440" *) reg2dp_kernel_height;
  assign _2340_ = bubble_add < (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) flush_in_next_surf;
  assign _1913_[2:0] = padding_stride_num * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1299" *) pooling_stride_v;
  assign pad_value = $signed(pad_table_out) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6289" *) $signed({ 1'b0, kernel_width_cfg });
  assign data_hmult_16bit_0_ext_ff = $signed(pout_data_0_0[21:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6366" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_hmult_16bit_1_ext_ff = $signed(pout_data_0_1[21:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6367" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_hmult_16bit_2_ext_ff = $signed(pout_data_0_2[21:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6368" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_hmult_16bit_3_ext_ff = $signed(pout_data_0_3[21:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6369" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_hmult_8bit_0_lsb_ext_ff = $signed(pout_data_0_0[13:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6571" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_hmult_8bit_0_msb_ext_ff = $signed(pout_data_0_0[27:14]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6572" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_hmult_8bit_1_lsb_ext_ff = $signed(pout_data_0_1[13:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6573" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_hmult_8bit_1_msb_ext_ff = $signed(pout_data_0_1[27:14]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6574" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_hmult_8bit_2_lsb_ext_ff = $signed(pout_data_0_2[13:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6575" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_hmult_8bit_2_msb_ext_ff = $signed(pout_data_0_2[27:14]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6576" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_hmult_8bit_3_lsb_ext_ff = $signed(pout_data_0_3[13:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6577" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_hmult_8bit_3_msb_ext_ff = $signed(pout_data_0_3[27:14]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6578" *) $signed({ 1'b0, reg2dp_recip_width_use });
  assign data_vmult_16bit_0_ext_ff = $signed(pout_data_stage0_0[18:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7021" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign data_vmult_16bit_1_ext_ff = $signed(pout_data_stage0_1[18:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7022" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign data_vmult_16bit_2_ext_ff = $signed(pout_data_stage0_2[18:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7023" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign data_vmult_16bit_3_ext_ff = $signed(pout_data_stage0_3[18:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7024" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign data_vmult_8bit_0_lsb_ext_ff = $signed(pout_data_stage0_0[10:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7226" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign data_vmult_8bit_0_msb_ext_ff = $signed(pout_data_stage0_0[21:11]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7227" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign data_vmult_8bit_1_lsb_ext_ff = $signed(pout_data_stage0_1[10:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7228" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign data_vmult_8bit_1_msb_ext_ff = $signed(pout_data_stage0_1[21:11]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7229" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign data_vmult_8bit_2_lsb_ext_ff = $signed(pout_data_stage0_2[10:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7230" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign data_vmult_8bit_2_msb_ext_ff = $signed(pout_data_stage0_2[21:11]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7231" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign data_vmult_8bit_3_lsb_ext_ff = $signed(pout_data_stage0_3[10:0]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7232" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign data_vmult_8bit_3_msb_ext_ff = $signed(pout_data_stage0_3[21:11]) * (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7233" *) $signed({ 1'b0, reg2dp_recip_height_use });
  assign splitw_enable = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1216" *) pooling_splitw_num_cfg;
  assign need_flush = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1493" *) flush_num;
  assign _2341_ = first_out_num != (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2166" *) 1'b1;
  assign _2342_ = pout_mem_size_v_use != (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6220" *) pooling_size_v_cfg;
  assign _2343_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1139" *) cur_datin_disable;
  assign _2344_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1140" *) one_width_disable;
  assign _2345_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1301" *) wr_total_cube_done;
  assign _2346_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1440" *) _3073_;
  assign _2347_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2076" *) is_one_width_in;
  assign _2348_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) cube_end_flag;
  assign _2349_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) need_bubble;
  assign _2350_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) wr_subcube_dat_done;
  assign _2351_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2332" *) last_pooling_flag;
  assign _2352_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2348" *) stride_trig_end;
  assign _2353_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0004_[15];
  assign _2354_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0005_[15];
  assign _2355_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0104_[15];
  assign _2356_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0105_[15];
  assign _2357_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0204_[15];
  assign _2358_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0205_[15];
  assign _2359_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0304_[15];
  assign _2360_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0305_[15];
  assign _2361_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0018_[15];
  assign _2362_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0118_[15];
  assign _2363_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0218_[15];
  assign _2364_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0318_[15];
  assign _2365_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0030_[15];
  assign _2366_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0130_[15];
  assign _2367_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0230_[15];
  assign _2368_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0330_[15];
  assign _2369_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0042_[15];
  assign _2370_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0142_[15];
  assign _2371_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0242_[15];
  assign _2372_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0342_[15];
  assign _2373_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0054_[15];
  assign _2374_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0154_[15];
  assign _2375_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0254_[15];
  assign _2376_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0354_[15];
  assign _2377_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0066_[15];
  assign _2378_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0166_[15];
  assign _2379_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0266_[15];
  assign _2380_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0366_[15];
  assign _2381_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0078_[15];
  assign _2382_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0178_[15];
  assign _2383_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0278_[15];
  assign _2384_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0378_[15];
  assign _2385_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0090_[15];
  assign _2386_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0190_[15];
  assign _2387_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0290_[15];
  assign _2388_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0390_[15];
  assign _2389_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) reg2dp_fp16_en;
  assign _2390_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0981_[0];
  assign _2391_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0984_[0];
  assign _2392_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0987_[0];
  assign _2393_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0990_[0];
  assign _2394_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0993_[0];
  assign _2395_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0996_[0];
  assign _2396_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0999_[0];
  assign _2397_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _1002_[0];
  assign _2398_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0981_[1];
  assign _2399_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0984_[1];
  assign _2400_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0987_[1];
  assign _2401_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0990_[1];
  assign _2402_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0993_[1];
  assign _2403_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0996_[1];
  assign _2404_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0999_[1];
  assign _2405_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _1002_[1];
  assign _2406_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0981_[2];
  assign _2407_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0984_[2];
  assign _2408_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0987_[2];
  assign _2409_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0990_[2];
  assign _2410_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0993_[2];
  assign _2411_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0996_[2];
  assign _2412_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0999_[2];
  assign _2413_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _1002_[2];
  assign _2414_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0981_[3];
  assign _2415_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0984_[3];
  assign _2416_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0987_[3];
  assign _2417_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0990_[3];
  assign _2418_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0993_[3];
  assign _2419_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0996_[3];
  assign _2420_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0999_[3];
  assign _2421_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _1002_[3];
  assign _2422_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4330" *) wr_data_stage0_vld;
  assign _2423_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4347" *) wr_data_stage1_vld;
  assign _2424_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4351" *) cur_datin_disable_d;
  assign _2425_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4351" *) one_width_disable_d;
  assign _2426_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4364" *) cur_datin_disable_2d;
  assign _2427_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4364" *) one_width_disable_2d;
  assign _2428_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4370" *) fp16_mean_pool_cfg;
  assign _2429_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4377" *) cur_datin_disable_3d;
  assign _2430_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4377" *) one_width_disable_3d;
  assign _2431_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5847" *) wr_data_stage2_vld;
  assign _2432_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5910" *) pout_data_stage1_vld;
  assign _2433_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5921" *) pout_data_stage2_vld;
  assign _2434_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5995" *) pout_data_stage3_vld;
  assign _2435_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6325" *) fp16_en;
  assign _2436_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6374" *) _3114_;
  assign _2437_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6374" *) data_hmult_16bit_0_ext[15];
  assign _2438_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6375" *) _3115_;
  assign _2439_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6375" *) data_hmult_16bit_1_ext[15];
  assign _2440_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6376" *) _3116_;
  assign _2441_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6376" *) data_hmult_16bit_2_ext[15];
  assign _2442_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6377" *) _3117_;
  assign _2443_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6377" *) data_hmult_16bit_3_ext[15];
  assign _2444_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6587" *) _3118_;
  assign _2445_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6587" *) data_hmult_8bit_0_lsb_ext[15];
  assign _2446_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6588" *) _3119_;
  assign _2447_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6588" *) data_hmult_8bit_0_msb_ext[15];
  assign _2448_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6589" *) _3120_;
  assign _2449_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6589" *) data_hmult_8bit_1_lsb_ext[15];
  assign _2450_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6590" *) _3121_;
  assign _2451_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6590" *) data_hmult_8bit_1_msb_ext[15];
  assign _2452_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6591" *) _3122_;
  assign _2453_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6591" *) data_hmult_8bit_2_lsb_ext[15];
  assign _2454_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6592" *) _3123_;
  assign _2455_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6592" *) data_hmult_8bit_2_msb_ext[15];
  assign _2456_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6593" *) _3124_;
  assign _2457_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6593" *) data_hmult_8bit_3_lsb_ext[15];
  assign _2458_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6594" *) _3125_;
  assign _2459_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6594" *) data_hmult_8bit_3_msb_ext[15];
  assign _2460_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7029" *) _3126_;
  assign _2461_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7029" *) data_vmult_16bit_0_ext[15];
  assign _2462_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7030" *) _3127_;
  assign _2463_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7030" *) data_vmult_16bit_1_ext[15];
  assign _2464_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7031" *) _3128_;
  assign _2465_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7031" *) data_vmult_16bit_2_ext[15];
  assign _2466_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7032" *) _3129_;
  assign _2467_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7032" *) data_vmult_16bit_3_ext[15];
  assign _2468_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7242" *) _3130_;
  assign _2469_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7242" *) data_vmult_8bit_0_lsb_ext[15];
  assign _2470_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7243" *) _3131_;
  assign _2471_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7243" *) data_vmult_8bit_0_msb_ext[15];
  assign _2472_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7244" *) _3132_;
  assign _2473_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7244" *) data_vmult_8bit_1_lsb_ext[15];
  assign _2474_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7245" *) _3133_;
  assign _2475_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7245" *) data_vmult_8bit_1_msb_ext[15];
  assign _2476_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7246" *) _3134_;
  assign _2477_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7246" *) data_vmult_8bit_2_lsb_ext[15];
  assign _2478_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7247" *) _3135_;
  assign _2479_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7247" *) data_vmult_8bit_2_msb_ext[15];
  assign _2480_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7248" *) _3136_;
  assign _2481_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7248" *) data_vmult_8bit_3_lsb_ext[15];
  assign _2482_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7249" *) _3137_;
  assign _2483_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7249" *) data_vmult_8bit_3_msb_ext[15];
  assign _2484_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7963" *) din_pd_d4[245];
  assign _2485_ = ~ (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7963" *) din_pd_d4[254];
  assign init_cnt = middle_surface_trig | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1303" *) pdp_op_start;
  assign _2486_ = init_cnt | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1325" *) stride_end;
  assign _2016_ = _2486_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1325" *) wr_line_dat_done;
  assign _2487_ = _2034_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) _2035_;
  assign _2488_ = _2487_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) _2036_;
  assign _2489_ = _2488_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) _2037_;
  assign _2490_ = _2489_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) _2038_;
  assign _2491_ = _2490_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) _2039_;
  assign _2492_ = _2040_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *) _2041_;
  assign _2493_ = _2492_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *) _2042_;
  assign _2494_ = _2493_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *) _2043_;
  assign _2495_ = _2494_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *) _2044_;
  assign _1929_[0] = _2495_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1776" *) _2045_;
  assign _2496_ = _2046_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) _2047_;
  assign _2497_ = _2496_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) _2048_;
  assign _2498_ = _2497_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) _2049_;
  assign _2499_ = _2498_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) _2050_;
  assign _2500_ = _2499_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) _2051_;
  assign _2501_ = _2052_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) _2053_;
  assign _2502_ = _2501_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) _2054_;
  assign _2503_ = _2502_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) _2055_;
  assign _2504_ = _2503_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) _2056_;
  assign _2505_ = _2504_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) _2057_;
  assign _2506_ = _2058_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *) _2059_;
  assign _2507_ = _2506_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *) _2060_;
  assign _2508_ = _2507_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *) _2061_;
  assign _2509_ = _2508_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *) _2062_;
  assign _1926_[0] = _2509_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1785" *) _2063_;
  assign _2510_ = _2064_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) _2065_;
  assign _2511_ = _2510_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) _2066_;
  assign _2512_ = _2511_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) _2067_;
  assign _2513_ = _2512_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) _2068_;
  assign _2514_ = _2513_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) _2069_;
  assign _2515_ = _2070_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) _2071_;
  assign _2516_ = _2515_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) _2072_;
  assign _2517_ = _2516_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) _2073_;
  assign _2518_ = _2517_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) _2074_;
  assign _2519_ = _2518_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) _2075_;
  assign _2520_ = _2076_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) _2077_;
  assign _2521_ = _2520_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) _2078_;
  assign _2522_ = _2521_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) _2079_;
  assign _2523_ = _2522_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) _2080_;
  assign _2524_ = _2523_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) _2081_;
  assign _2525_ = _2082_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *) _2083_;
  assign _2526_ = _2525_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *) _2084_;
  assign _2527_ = _2526_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *) _2085_;
  assign _2528_ = _2527_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *) _2086_;
  assign _1923_[0] = _2528_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1796" *) _2087_;
  assign _2529_ = _2088_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) _2089_;
  assign _2530_ = _2529_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) _2090_;
  assign _2531_ = _2530_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) _2091_;
  assign _2532_ = _2531_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) _2092_;
  assign _2533_ = _2532_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) _2093_;
  assign _2534_ = _2094_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) _2095_;
  assign _2535_ = _2534_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) _2096_;
  assign _2536_ = _2535_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) _2097_;
  assign _2537_ = _2536_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) _2098_;
  assign _2538_ = _2537_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) _2099_;
  assign _2539_ = _2100_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) _2101_;
  assign _2540_ = _2539_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) _2102_;
  assign _2541_ = _2540_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) _2103_;
  assign _2542_ = _2541_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) _2104_;
  assign _2543_ = _2542_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) _2105_;
  assign _2544_ = _2106_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) _2107_;
  assign _2545_ = _2544_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) _2108_;
  assign _2546_ = _2545_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) _2109_;
  assign _2547_ = _2546_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) _2110_;
  assign _2548_ = _2547_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) _2111_;
  assign _2549_ = _2112_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *) _2113_;
  assign _2550_ = _2549_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *) _2114_;
  assign _2551_ = _2550_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *) _2115_;
  assign _2552_ = _2551_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *) _2116_;
  assign _1920_[0] = _2552_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1809" *) _2117_;
  assign _2553_ = _2118_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) _2119_;
  assign _2554_ = _2553_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) _2120_;
  assign _2555_ = _2554_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) _2121_;
  assign _2556_ = _2555_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) _2122_;
  assign _2557_ = _2556_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) _2123_;
  assign _2558_ = _2124_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) _2125_;
  assign _2559_ = _2558_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) _2126_;
  assign _2560_ = _2559_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) _2127_;
  assign _2561_ = _2560_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) _2128_;
  assign _2562_ = _2561_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) _2129_;
  assign _2563_ = _2130_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) _2131_;
  assign _2564_ = _2563_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) _2132_;
  assign _2565_ = _2564_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) _2133_;
  assign _2566_ = _2565_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) _2134_;
  assign _2567_ = _2566_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) _2135_;
  assign _2568_ = _2136_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) _2137_;
  assign _2569_ = _2568_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) _2138_;
  assign _2570_ = _2569_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) _2139_;
  assign _2571_ = _2570_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) _2140_;
  assign _2572_ = _2571_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) _2141_;
  assign _2573_ = _2142_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) _2143_;
  assign _2574_ = _2573_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) _2144_;
  assign _2575_ = _2574_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) _2145_;
  assign _2576_ = _2575_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) _2146_;
  assign _2577_ = _2576_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) _2147_;
  assign _2578_ = _2148_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *) _2149_;
  assign _2579_ = _2578_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *) _2150_;
  assign _2580_ = _2579_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *) _2151_;
  assign _2581_ = _2580_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *) _2152_;
  assign _1917_[0] = _2581_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1824" *) _2153_;
  assign _2582_ = _2154_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) _2155_;
  assign _2583_ = _2582_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) _2156_;
  assign _2584_ = _2583_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) _2157_;
  assign _2585_ = _2584_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) _2158_;
  assign _2586_ = _2585_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) _2159_;
  assign _2587_ = _2160_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) _2161_;
  assign _2588_ = _2587_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) _2162_;
  assign _2589_ = _2588_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) _2163_;
  assign _2590_ = _2589_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) _2164_;
  assign _2591_ = _2590_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) _2165_;
  assign _2592_ = _2166_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) _2167_;
  assign _2593_ = _2592_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) _2168_;
  assign _2594_ = _2593_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) _2169_;
  assign _2595_ = _2594_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) _2170_;
  assign _2596_ = _2595_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) _2171_;
  assign _2597_ = _2172_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) _2173_;
  assign _2598_ = _2597_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) _2174_;
  assign _2599_ = _2598_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) _2175_;
  assign _2600_ = _2599_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) _2176_;
  assign _2601_ = _2600_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) _2177_;
  assign _2602_ = _2178_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) _2179_;
  assign _2603_ = _2602_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) _2180_;
  assign _2604_ = _2603_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) _2181_;
  assign _2605_ = _2604_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) _2182_;
  assign _2606_ = _2605_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) _2183_;
  assign _2607_ = _2184_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) _2185_;
  assign _2608_ = _2607_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) _2186_;
  assign _2609_ = _2608_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) _2187_;
  assign _2610_ = _2609_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) _2188_;
  assign _2611_ = _2610_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) _2189_;
  assign _2612_ = _2190_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *) _2191_;
  assign _2613_ = _2612_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *) _2192_;
  assign _2614_ = _2613_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *) _2193_;
  assign _2615_ = _2614_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *) _2194_;
  assign _1914_[0] = _2615_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1841" *) _2195_;
  assign _2616_ = _2207_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1981" *) _2209_;
  assign _2617_ = _2209_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2007" *) _2211_;
  assign _2618_ = _2617_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2033" *) _2213_;
  assign _2619_ = _1293_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2076" *) _1294_;
  assign _2620_ = _1295_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2078" *) _1296_;
  assign _2621_ = _1299_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) _1302_;
  assign _2622_ = _1303_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2182" *) _1304_;
  assign _2623_ = pooling_2d_rdy | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2313" *) wr_surface_dat_done;
  assign unit2d_set[0] = unit2d_set_trig[0] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2333" *) init_unit2d_set[0];
  assign unit2d_clr[0] = _1308_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2334" *) wr_surface_dat_done;
  assign unit2d_set[1] = unit2d_set_trig[1] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2349" *) init_unit2d_set[1];
  assign unit2d_clr[1] = _1311_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2350" *) wr_surface_dat_done;
  assign unit2d_set[2] = unit2d_set_trig[2] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2365" *) init_unit2d_set[2];
  assign unit2d_clr[2] = _1314_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2366" *) wr_surface_dat_done;
  assign unit2d_set[3] = unit2d_set_trig[3] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2381" *) init_unit2d_set[3];
  assign unit2d_clr[3] = _1317_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2382" *) wr_surface_dat_done;
  assign unit2d_set[4] = unit2d_set_trig[4] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2397" *) init_unit2d_set[4];
  assign unit2d_clr[4] = _1320_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2398" *) wr_surface_dat_done;
  assign unit2d_set[5] = unit2d_set_trig[5] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2413" *) init_unit2d_set[5];
  assign unit2d_clr[5] = _1323_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2414" *) wr_surface_dat_done;
  assign unit2d_set[6] = unit2d_set_trig[6] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2429" *) init_unit2d_set[6];
  assign unit2d_clr[6] = _1326_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2430" *) wr_surface_dat_done;
  assign unit2d_set[7] = unit2d_set_trig[7] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2445" *) init_unit2d_set[7];
  assign unit2d_clr[7] = _1329_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2446" *) wr_surface_dat_done;
  assign _2624_ = unit2d_vsize1_0 | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2764" *) unit2d_vsize2_0;
  assign _2625_ = _2624_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2764" *) unit2d_vsize3_0;
  assign unit2d_vsize_0 = _2625_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2764" *) unit2d_vsize4_0;
  assign unit2d_vsize_1 = _2625_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2765" *) unit2d_vsize4_1;
  assign _2626_ = _2624_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2766" *) unit2d_vsize3_2;
  assign unit2d_vsize_2 = _2626_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2766" *) unit2d_vsize4_2;
  assign unit2d_vsize_3 = _2626_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2767" *) unit2d_vsize4_3;
  assign _2627_ = unit2d_vsize1_0 | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2768" *) unit2d_vsize2_4;
  assign _2628_ = _2627_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2768" *) unit2d_vsize3_4;
  assign unit2d_vsize_4 = _2628_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2768" *) unit2d_vsize4_4;
  assign unit2d_vsize_5 = _2628_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2769" *) unit2d_vsize4_5;
  assign _2629_ = _2627_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2770" *) unit2d_vsize3_6;
  assign unit2d_vsize_6 = _2629_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2770" *) unit2d_vsize4_6;
  assign unit2d_vsize_7 = _2629_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2771" *) unit2d_vsize4_7;
  assign active_last_line = _2224_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3261" *) last_line_in;
  assign _1054_ = _2248_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3405" *) _2249_;
  assign _2630_ = mem_re1 | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3412" *) mem_re2;
  assign _2631_ = _2630_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3412" *) mem_re3;
  assign mem_re = _2631_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3412" *) mem_re4;
  assign _2632_ = { mem_re1_1st[7], mem_re1_1st[7], mem_re1_1st[7], mem_re1_1st[7], mem_re1_1st[7], mem_re1_1st[7], mem_re1_1st[7], mem_re1_1st[7] } | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3413" *) { mem_re2_1st[7], mem_re2_1st[7], mem_re2_1st[7], mem_re2_1st[7], mem_re2_1st[3], mem_re2_1st[3], mem_re2_1st[3], mem_re2_1st[3] };
  assign _2633_ = _2632_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3413" *) { mem_re3_1st[7], mem_re3_1st[7], mem_re3_1st[5], mem_re3_1st[5], mem_re3_1st[3], mem_re3_1st[3], mem_re3_1st[1], mem_re3_1st[1] };
  assign mem_re_1st = _2633_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3413" *) mem_re4_1st;
  assign _2634_ = wr_line_dat_done | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3420" *) last_sub_lbuf_done;
  assign _2635_ = _2634_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3420" *) line_end;
  assign _2636_ = sub_lbuf_dout_done | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3432" *) wr_line_dat_done;
  assign _2637_ = _2636_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3432" *) line_end;
  assign _2262_ = load_din | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3435" *) _1366_;
  assign _0981_ = _0977_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3594" *) _0978_;
  assign _0984_ = _0977_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3594" *) _0983_;
  assign _0987_ = _0977_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3594" *) _0986_;
  assign _0990_ = _0977_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3594" *) _0989_;
  assign _0993_ = _0977_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3594" *) _0992_;
  assign _0996_ = _0977_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3594" *) _0995_;
  assign _0999_ = _0977_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3594" *) _0998_;
  assign _1002_ = _0977_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3594" *) _1001_;
  assign _2638_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _1671_;
  assign _2639_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _1672_;
  assign _2640_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _1673_;
  assign _2641_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _1674_;
  assign _2642_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _1675_;
  assign _2643_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _1676_;
  assign _2644_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _1677_;
  assign _2645_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _1678_;
  assign _2646_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _1679_;
  assign _2647_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _1680_;
  assign _2648_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _1681_;
  assign _2649_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _1682_;
  assign _2650_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _1683_;
  assign _2651_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _1684_;
  assign _2652_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _1685_;
  assign _2653_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _1686_;
  assign _2654_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _1687_;
  assign _2655_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _1688_;
  assign _2656_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _1689_;
  assign _2657_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _1690_;
  assign _2658_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _1691_;
  assign _2659_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _1692_;
  assign _2660_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _1693_;
  assign _2661_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _1694_;
  assign _2662_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _1695_;
  assign _2663_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _1696_;
  assign _2664_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _1697_;
  assign _2665_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _1698_;
  assign _2666_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _1699_;
  assign _2667_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _1700_;
  assign _2668_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _1701_;
  assign _2669_ = _2389_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _1702_;
  assign _2252_ = _3110_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4148" *) _1704_;
  assign pooling1d_norm_rdy = _2422_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4330" *) wr_data_stage0_prdy;
  assign _2670_ = one_width_disable | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4333" *) cur_datin_disable;
  assign wr_data_stage0_prdy = _2423_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4347" *) wr_data_stage1_prdy;
  assign _2671_ = mem_re[0] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4582" *) mem_re_last[0];
  assign _2672_ = mem_re[1] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4592" *) mem_re_last[1];
  assign _2673_ = mem_re[2] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4602" *) mem_re_last[2];
  assign _2674_ = mem_re[3] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4612" *) mem_re_last[3];
  assign _2675_ = mem_re[4] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4622" *) mem_re_last[4];
  assign _2676_ = mem_re[5] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4632" *) mem_re_last[5];
  assign _2677_ = mem_re[6] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4642" *) mem_re_last[6];
  assign _2678_ = mem_re[7] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4652" *) mem_re_last[7];
  assign _2679_ = _1710_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5041" *) _1711_;
  assign _2680_ = cur_datin_disable | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5052" *) last_out_en;
  assign _2681_ = mem_re2_last | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5085" *) mem_re3_last;
  assign mem_re_last = _2681_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5085" *) mem_re4_last;
  assign _2261_ = _1729_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5090" *) _1366_;
  assign _2263_ = load_wr_stage1 | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5395" *) _1730_;
  assign _2264_ = _1731_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5456" *) _1730_;
  assign _2682_ = load_wr_stage2 | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5764" *) _1732_;
  assign _2683_ = pout_mem_data_sel_3_last | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5790" *) pout_mem_data_sel_2_last;
  assign pout_mem_data_sel_last = _2683_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5790" *) pout_mem_data_sel_1_last;
  assign _2684_ = _1762_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5792" *) _1763_;
  assign _2685_ = _2684_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5793" *) _1764_;
  assign _2686_ = _2685_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5794" *) _1765_;
  assign _2687_ = _2686_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5795" *) _1766_;
  assign _2688_ = _2687_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5796" *) _1767_;
  assign _2689_ = _2688_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5797" *) _1768_;
  assign pout_mem_data_last = _2689_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5798" *) _1769_;
  assign _2690_ = rd_line_out_done | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5810" *) rd_sub_lbuf_end;
  assign rd_sub_lbuf_end = _1770_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5816" *) rd_line_out_done;
  assign rd_comb_lbuf_end = _1771_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5828" *) rd_line_out_done;
  assign _2691_ = rd_lbuf_end | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5835" *) _1772_;
  assign _2692_ = _1775_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5845" *) _1732_;
  assign rd_pout_data_en = rd_line_out | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5845" *) _2692_;
  assign _2693_ = _2431_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5847" *) pout_data_stage0_prdy;
  assign pout_data_stage0_prdy = _2432_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5910" *) pout_data_stage1_prdy;
  assign pout_data_stage1_prdy = _2433_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5921" *) pout_data_stage2_prdy;
  assign pout_data_stage2_prdy = _2434_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5995" *) pout_data_stage3_prdy;
  assign _2694_ = pout_mem_data_sel_3 | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6160" *) pout_mem_data_sel_2;
  assign _2695_ = _2694_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6160" *) pout_mem_data_sel_1;
  assign pout_mem_data_sel = _2695_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6160" *) pout_mem_data_sel_0;
  assign int_pout_mem_data = pout_mem_data_act | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6192" *) pout_mem_data_last;
  assign _2696_ = _1829_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6374" *) _2437_;
  assign _2697_ = _1830_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6375" *) _2439_;
  assign _2698_ = _1831_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6376" *) _2441_;
  assign _2699_ = _1832_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6377" *) _2443_;
  assign _2700_ = _1837_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6587" *) _2445_;
  assign _2701_ = _1838_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6588" *) _2447_;
  assign _2702_ = _1839_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6589" *) _2449_;
  assign _2703_ = _1840_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6590" *) _2451_;
  assign _2704_ = _1841_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6591" *) _2453_;
  assign _2705_ = _1842_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6592" *) _2455_;
  assign _2706_ = _1843_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6593" *) _2457_;
  assign _2707_ = _1844_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6594" *) _2459_;
  assign _2708_ = _1853_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7029" *) _2461_;
  assign _2709_ = _1854_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7030" *) _2463_;
  assign _2710_ = _1855_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7031" *) _2465_;
  assign _2711_ = _1856_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7032" *) _2467_;
  assign _2712_ = _1861_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7242" *) _2469_;
  assign _2713_ = _1862_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7243" *) _2471_;
  assign _2714_ = _1863_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7244" *) _2473_;
  assign _2715_ = _1864_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7245" *) _2475_;
  assign _2716_ = _1865_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7246" *) _2477_;
  assign _2717_ = _1866_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7247" *) _2479_;
  assign _2718_ = _1867_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7248" *) _2481_;
  assign _2719_ = _1868_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7249" *) _2483_;
  assign _2720_ = _3525_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8025" *) _3526_;
  assign _2721_ = _2720_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8026" *) _3527_;
  assign _2722_ = _2721_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8027" *) _3528_;
  assign _2723_ = _2722_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8028" *) _3529_;
  assign _2724_ = _2723_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8029" *) _3530_;
  assign _2725_ = _2724_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8030" *) _3531_;
  assign fp_pout_mem_data_act = _2725_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8030" *) _3532_;
  assign _2726_ = _3533_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8033" *) _3534_;
  assign _2727_ = _2726_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8034" *) _3535_;
  assign _2728_ = _2727_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8035" *) _3536_;
  assign _2729_ = _2728_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8036" *) _3537_;
  assign _2730_ = _2729_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8037" *) _3538_;
  assign _2731_ = _2730_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8038" *) _3539_;
  assign fp_pout_mem_data_last = _2731_ | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8038" *) _3540_;
  assign fp16_mul_pad_line_in_pd_d0 = fp_pout_mem_data_act | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8039" *) fp_pout_mem_data_last;
  assign _2732_ = din_pd_d4[128:121] | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8762" *) din_pd_d4[168:161];
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_stage1_0 <= 16'b0000000000000000;
    else
      pout_data_stage1_0 <= _1085_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_stage1_1 <= 16'b0000000000000000;
    else
      pout_data_stage1_1 <= _1086_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_stage1_2 <= 16'b0000000000000000;
    else
      pout_data_stage1_2 <= _1087_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_stage1_3 <= 16'b0000000000000000;
    else
      pout_data_stage1_3 <= _1088_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_stage0_0 <= 22'b0000000000000000000000;
    else
      pout_data_stage0_0 <= _1081_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_stage0_1 <= 22'b0000000000000000000000;
    else
      pout_data_stage0_1 <= _1082_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_stage0_2 <= 22'b0000000000000000000000;
    else
      pout_data_stage0_2 <= _1083_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_stage0_3 <= 22'b0000000000000000000000;
    else
      pout_data_stage0_3 <= _1084_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg2dp_recip_height_use <= 17'b00000000000000000;
    else
      reg2dp_recip_height_use <= reg2dp_recip_height_cfg;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      reg2dp_recip_width_use <= 17'b00000000000000000;
    else
      reg2dp_recip_width_use <= reg2dp_recip_width_cfg;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_0_0 <= 28'b0000000000000000000000000000;
    else
      pout_data_0_0 <= _1077_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_0_1 <= 28'b0000000000000000000000000000;
    else
      pout_data_0_1 <= _1078_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_0_2 <= 28'b0000000000000000000000000000;
    else
      pout_data_0_2 <= _1079_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_0_3 <= 28'b0000000000000000000000000000;
    else
      pout_data_0_3 <= _1080_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_mem_data_0 <= 28'b0000000000000000000000000000;
    else
      pout_mem_data_0 <= _1092_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_mem_data_1 <= 28'b0000000000000000000000000000;
    else
      pout_mem_data_1 <= _1093_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_mem_data_2 <= 28'b0000000000000000000000000000;
    else
      pout_mem_data_2 <= _1094_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_mem_data_3 <= 28'b0000000000000000000000000000;
    else
      pout_mem_data_3 <= _1095_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_mem_size_v <= 3'b000;
    else
      pout_mem_size_v <= _1096_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_stage3_vld <= 1'b0;
    else
      pout_data_stage3_vld <= _1091_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_pout_data_en_4d <= 1'b0;
    else
      rd_pout_data_en_4d <= _1102_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_pout_data_en_3d <= 1'b0;
    else
      rd_pout_data_en_3d <= _1101_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_stage2_vld <= 1'b0;
    else
      pout_data_stage2_vld <= _1090_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_pout_data_en_2d <= 1'b0;
    else
      rd_pout_data_en_2d <= _1100_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_data_stage1_vld <= 1'b0;
    else
      pout_data_stage1_vld <= _1089_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_pout_data_en_d <= 1'b0;
    else
      rd_pout_data_en_d <= _1103_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_comb_lbuf_cnt <= 3'b000;
    else
      rd_comb_lbuf_cnt <= _1098_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_sub_lbuf_cnt <= 3'b000;
    else
      rd_sub_lbuf_cnt <= _1104_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_line_out_cnt <= 6'b000000;
    else
      rd_line_out_cnt <= _1099_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      one_width_disable_3d <= 1'b0;
    else
      one_width_disable_3d <= _1068_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cur_datin_disable_3d <= 1'b0;
    else
      cur_datin_disable_3d <= _1013_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      one_width_disable_2d <= 1'b0;
    else
      one_width_disable_2d <= _1067_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cur_datin_disable_2d <= 1'b0;
    else
      cur_datin_disable_2d <= _1012_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_cnt_pooling_last_2d <= 3'b000;
    else
      unit2d_cnt_pooling_last_2d <= _1113_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re_last_2d <= 8'b00000000;
    else
      mem_re_last_2d <= _1062_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      one_width_disable_d <= 1'b0;
    else
      one_width_disable_d <= _1069_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cur_datin_disable_d <= 1'b0;
    else
      cur_datin_disable_d <= _1014_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_cnt_pooling_last_d <= 3'b000;
    else
      unit2d_cnt_pooling_last_d <= _1114_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re_last_d <= 8'b00000000;
    else
      mem_re_last_d <= _1063_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      flush_read_en_d <= 1'b0;
    else
      flush_read_en_d <= _1017_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re2_sel_last <= 1'b0;
    else
      mem_re2_sel_last <= _1053_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re3_sel_last <= 1'b0;
    else
      mem_re3_sel_last <= _1055_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re4_sel_last <= 1'b0;
    else
      mem_re4_sel_last <= _1057_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_cnt_pooling_last <= 3'b000;
    else
      unit2d_cnt_pooling_last <= _1112_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      int_mem_waddr <= 6'b000000;
    else
      int_mem_waddr <= _1018_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      int_mem_we <= 8'b00000000;
    else
      int_mem_we <= _1027_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      int_mem_wdata_0 <= 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      int_mem_wdata_0 <= _1019_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      int_mem_wdata_1 <= 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      int_mem_wdata_1 <= _1020_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      int_mem_wdata_2 <= 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      int_mem_wdata_2 <= _1021_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      int_mem_wdata_3 <= 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      int_mem_wdata_3 <= _1022_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      int_mem_wdata_4 <= 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      int_mem_wdata_4 <= _1023_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      int_mem_wdata_5 <= 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      int_mem_wdata_5 <= _1024_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      int_mem_wdata_6 <= 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      int_mem_wdata_6 <= _1025_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      int_mem_wdata_7 <= 116'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      int_mem_wdata_7 <= _1026_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wr_data_stage2_vld <= 1'b0;
    else
      wr_data_stage2_vld <= _1155_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wr_data_stage1_vld <= 1'b0;
    else
      wr_data_stage1_vld <= _1154_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wr_data_stage0_vld <= 1'b0;
    else
      wr_data_stage0_vld <= _1153_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re_2d <= 8'b00000000;
    else
      mem_re_2d <= _1060_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re_d <= 8'b00000000;
    else
      mem_re_d <= _1061_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_raddr_d <= 6'b000000;
    else
      mem_raddr_d <= _1050_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re_1st_2d <= 8'b00000000;
    else
      mem_re_1st_2d <= _1058_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re_1st_d <= 8'b00000000;
    else
      mem_re_1st_d <= _1059_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      last_active_line_2d <= 1'b0;
    else
      last_active_line_2d <= _1028_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      last_active_line_d <= 1'b0;
    else
      last_active_line_d <= _1029_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wr_surface_dat_done_2d <= 1'b0;
    else
      wr_surface_dat_done_2d <= _1162_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_raddr_2d <= 6'b000000;
    else
      mem_raddr_2d <= _1049_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wr_line_end_2d <= 1'b0;
    else
      wr_line_end_2d <= _1157_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      datin_buf_2d <= 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      datin_buf_2d <= _1016_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data0 <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data0 <= _1033_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data1 <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data1 <= _1035_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data2 <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data2 <= _1037_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data3 <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data3 <= _1039_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data4 <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data4 <= _1041_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data5 <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data5 <= _1043_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data6 <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data6 <= _1045_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data7 <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data7 <= _1047_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data0_lst <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data0_lst <= _1034_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data1_lst <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data1_lst <= _1036_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data2_lst <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data2_lst <= _1038_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data3_lst <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data3_lst <= _1040_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data4_lst <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data4_lst <= _1042_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data5_lst <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data5_lst <= _1044_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data6_lst <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data6_lst <= _1046_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_data7_lst <= 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      mem_data7_lst <= _1048_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sub_lbuf_dout_cnt <= 6'b000000;
    else
      sub_lbuf_dout_cnt <= _1107_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wr_sub_lbuf_cnt <= 3'b000;
    else
      wr_sub_lbuf_cnt <= _1160_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re1_sel <= 1'b0;
    else
      mem_re1_sel <= _1051_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re2_sel <= 1'b0;
    else
      mem_re2_sel <= _1052_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re3_sel <= 1'b0;
    else
      mem_re3_sel <= _1054_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      mem_re4_sel <= 1'b0;
    else
      mem_re4_sel <= _1056_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_mem_1strd[7] <= 1'b0;
    else
      unit2d_mem_1strd[7] <= _1131_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_mem_1strd[6] <= 1'b0;
    else
      unit2d_mem_1strd[6] <= _1130_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_mem_1strd[5] <= 1'b0;
    else
      unit2d_mem_1strd[5] <= _1129_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_mem_1strd[4] <= 1'b0;
    else
      unit2d_mem_1strd[4] <= _1128_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_mem_1strd[3] <= 1'b0;
    else
      unit2d_mem_1strd[3] <= _1127_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_mem_1strd[2] <= 1'b0;
    else
      unit2d_mem_1strd[2] <= _1126_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_mem_1strd[1] <= 1'b0;
    else
      unit2d_mem_1strd[1] <= _1125_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_mem_1strd[0] <= 1'b0;
    else
      unit2d_mem_1strd[0] <= _1124_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_7_d <= 3'b000;
    else
      unit2d_vsize_cnt_7_d <= _1147_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_6_d <= 3'b000;
    else
      unit2d_vsize_cnt_6_d <= _1145_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_5_d <= 3'b000;
    else
      unit2d_vsize_cnt_5_d <= _1143_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_4_d <= 3'b000;
    else
      unit2d_vsize_cnt_4_d <= _1141_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_3_d <= 3'b000;
    else
      unit2d_vsize_cnt_3_d <= _1139_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_2_d <= 3'b000;
    else
      unit2d_vsize_cnt_2_d <= _1137_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_1_d <= 3'b000;
    else
      unit2d_vsize_cnt_1_d <= _1135_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_0_d <= 3'b000;
    else
      unit2d_vsize_cnt_0_d <= _1133_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_7 <= 3'b000;
    else
      unit2d_vsize_cnt_7 <= _1146_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_6 <= 3'b000;
    else
      unit2d_vsize_cnt_6 <= _1144_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_5 <= 3'b000;
    else
      unit2d_vsize_cnt_5 <= _1142_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_4 <= 3'b000;
    else
      unit2d_vsize_cnt_4 <= _1140_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_3 <= 3'b000;
    else
      unit2d_vsize_cnt_3 <= _1138_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_2 <= 3'b000;
    else
      unit2d_vsize_cnt_2 <= _1136_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_1 <= 3'b000;
    else
      unit2d_vsize_cnt_1 <= _1134_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_vsize_cnt_0 <= 3'b000;
    else
      unit2d_vsize_cnt_0 <= _1132_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wr_surface_dat_done_buf <= 1'b0;
    else
      wr_surface_dat_done_buf <= _1163_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wr_line_end_buf <= 1'b0;
    else
      wr_line_end_buf <= _1158_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      datin_buf <= 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      datin_buf <= _1015_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_en[7] <= 1'b0;
    else
      unit2d_en[7] <= _1123_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_en[6] <= 1'b0;
    else
      unit2d_en[6] <= _1122_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_en[5] <= 1'b0;
    else
      unit2d_en[5] <= _1121_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_en[4] <= 1'b0;
    else
      unit2d_en[4] <= _1120_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_en[3] <= 1'b0;
    else
      unit2d_en[3] <= _1119_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_en[2] <= 1'b0;
    else
      unit2d_en[2] <= _1118_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_en[1] <= 1'b0;
    else
      unit2d_en[1] <= _1117_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_en[0] <= 1'b0;
    else
      unit2d_en[0] <= _1116_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_cnt_pooling <= 3'b000;
    else
      unit2d_cnt_pooling <= _1111_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      unit2d_cnt_stride <= 3'b000;
    else
      unit2d_cnt_stride <= _1115_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      one_width_bubble_cnt <= 3'b000;
    else
      one_width_bubble_cnt <= _1065_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      one_width_disable <= 1'b0;
    else
      one_width_disable <= _1066_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      last_out_cnt <= 3'b000;
    else
      last_out_cnt <= _1030_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      last_out_en <= 1'b0;
    else
      last_out_en <= _1031_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cube_end_flag <= 1'b0;
    else
      cube_end_flag <= _1010_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      bubble_cnt <= 3'b000;
    else
      bubble_cnt <= _1004_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      line_cnt <= 13'b0000000000000;
    else
      line_cnt <= _1032_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      channel_cnt <= 2'b00;
    else
      channel_cnt <= _1009_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      pout_width_cur_latch <= 13'b0000000000000;
    else
      pout_width_cur_latch <= _1097_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cur_datin_disable <= 1'b0;
    else
      cur_datin_disable <= _1011_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      surfend_need_bubble_flg <= 1'b0;
    else
      surfend_need_bubble_flg <= _1110_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      subend_need_flush_flg <= 1'b0;
    else
      subend_need_flush_flg <= _1108_;
  always @(posedge nvdla_core_clk)
      up_pnum1 <= _1148_;
  always @(posedge nvdla_core_clk)
      up_pnum2 <= _1149_;
  always @(posedge nvdla_core_clk)
      up_pnum3 <= _1150_;
  always @(posedge nvdla_core_clk)
      up_pnum4 <= _1151_;
  always @(posedge nvdla_core_clk)
      up_pnum5 <= _1152_;
  always @(posedge nvdla_core_clk)
      pnum_flush0 <= _1070_;
  always @(posedge nvdla_core_clk)
      pnum_flush1 <= _1071_;
  always @(posedge nvdla_core_clk)
      pnum_flush2 <= _1072_;
  always @(posedge nvdla_core_clk)
      pnum_flush3 <= _1073_;
  always @(posedge nvdla_core_clk)
      pnum_flush4 <= _1074_;
  always @(posedge nvdla_core_clk)
      pnum_flush5 <= _1075_;
  always @(posedge nvdla_core_clk)
      pnum_flush6 <= _1076_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      bubble_add <= 3'b000;
    else
      bubble_add <= _1003_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      bubble_num <= 3'b000;
    else
      bubble_num <= _1005_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      need_bubble <= 1'b0;
    else
      need_bubble <= _1064_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      bubble_num_use <= 3'b000;
    else
      bubble_num_use <= _1006_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      strip_ycnt_psize <= 3'b000;
    else
      strip_ycnt_psize <= _1105_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      strip_ycnt_stride <= 4'b0000;
    else
      strip_ycnt_stride <= _1106_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      buffer_lines_num <= 4'b0000;
    else
      buffer_lines_num <= _1007_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wr_splitc_cnt <= 8'b00000000;
    else
      wr_splitc_cnt <= _1159_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      surface_cnt_rd <= 11'b00000000000;
    else
      surface_cnt_rd <= _1109_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wr_surface_dat_cnt <= 13'b0000000000000;
    else
      wr_surface_dat_cnt <= _1161_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      wr_line_dat_cnt <= 13'b0000000000000;
    else
      wr_line_dat_cnt <= _1156_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      c_cnt <= 2'b00;
    else
      c_cnt <= _1008_;
  function [16:0] _5900_;
    input [16:0] a;
    input [118:0] b;
    input [6:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8780|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8772" *)
    (* parallel_case *)
    casez (s)
      7'b??????1:
        _5900_ = b[16:0];
      7'b?????1?:
        _5900_ = b[33:17];
      7'b????1??:
        _5900_ = b[50:34];
      7'b???1???:
        _5900_ = b[67:51];
      7'b??1????:
        _5900_ = b[84:68];
      7'b?1?????:
        _5900_ = b[101:85];
      7'b1??????:
        _5900_ = b[118:102];
      default:
        _5900_ = a;
    endcase
  endfunction
  assign kernel_width_fp17 = _5900_(17'b00111110000000000, 119'b01000000000000000010000010000000000100001000000000001000010100000000010000110000000000100001110000000001000100000000000, { _2739_, _2738_, _2737_, _2736_, _2735_, _2734_, _2733_ });
  assign _2733_ = reg2dp_kernel_width == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8780|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8772" *) 3'b111;
  assign _2734_ = reg2dp_kernel_width == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8779|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8772" *) 3'b110;
  assign _2735_ = reg2dp_kernel_width == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8778|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8772" *) 3'b101;
  assign _2736_ = reg2dp_kernel_width == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8777|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8772" *) 3'b100;
  assign _2737_ = reg2dp_kernel_width == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8776|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8772" *) 2'b11;
  assign _2738_ = reg2dp_kernel_width == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8775|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8772" *) 2'b10;
  assign _2739_ = reg2dp_kernel_width == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8774|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8772" *) 1'b1;
  assign _2740_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7657" *) { pout_data_stage0_3[18:11], pout_data_stage0_3[7:0] } : pout_data_stage0_3[15:0];
  assign _2741_ = rd_pout_data_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7656" *) _2740_ : pout_data_stage1_3;
  assign _2742_ = rd_pout_data_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7650" *) data_mult_stage1_in3 : pout_data_stage1_3;
  assign _1088_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7649" *) _2742_ : _2741_;
  assign _2743_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7657" *) { pout_data_stage0_2[18:11], pout_data_stage0_2[7:0] } : pout_data_stage0_2[15:0];
  assign _2744_ = rd_pout_data_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7656" *) _2743_ : pout_data_stage1_2;
  assign _2745_ = rd_pout_data_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7650" *) data_mult_stage1_in2 : pout_data_stage1_2;
  assign _1087_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7649" *) _2745_ : _2744_;
  assign _2746_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7657" *) { pout_data_stage0_1[18:11], pout_data_stage0_1[7:0] } : pout_data_stage0_1[15:0];
  assign _2747_ = rd_pout_data_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7656" *) _2746_ : pout_data_stage1_1;
  assign _2748_ = rd_pout_data_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7650" *) data_mult_stage1_in1 : pout_data_stage1_1;
  assign _1086_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7649" *) _2748_ : _2747_;
  assign _2749_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7657" *) { pout_data_stage0_0[18:11], pout_data_stage0_0[7:0] } : pout_data_stage0_0[15:0];
  assign _2750_ = rd_pout_data_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7656" *) _2749_ : pout_data_stage1_0;
  assign _2751_ = rd_pout_data_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7650" *) data_mult_stage1_in0 : pout_data_stage1_0;
  assign _1085_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7649" *) _2751_ : _2750_;
  assign _2752_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7004" *) { pout_data_0_3[24:14], pout_data_0_3[10:0] } : pout_data_0_3[21:0];
  assign _2753_ = rd_pout_data_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7003" *) _2752_ : pout_data_stage0_3;
  assign _2754_ = rd_pout_data_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6997" *) data_hmult_stage0_in3 : pout_data_stage0_3;
  assign _1084_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6996" *) _2754_ : _2753_;
  assign _2755_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7004" *) { pout_data_0_2[24:14], pout_data_0_2[10:0] } : pout_data_0_2[21:0];
  assign _2756_ = rd_pout_data_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7003" *) _2755_ : pout_data_stage0_2;
  assign _2757_ = rd_pout_data_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6997" *) data_hmult_stage0_in2 : pout_data_stage0_2;
  assign _1083_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6996" *) _2757_ : _2756_;
  assign _2758_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7004" *) { pout_data_0_1[24:14], pout_data_0_1[10:0] } : pout_data_0_1[21:0];
  assign _2759_ = rd_pout_data_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7003" *) _2758_ : pout_data_stage0_1;
  assign _2760_ = rd_pout_data_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6997" *) data_hmult_stage0_in1 : pout_data_stage0_1;
  assign _1082_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6996" *) _2760_ : _2759_;
  assign _2761_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7004" *) { pout_data_0_0[24:14], pout_data_0_0[10:0] } : pout_data_0_0[21:0];
  assign _2762_ = rd_pout_data_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7003" *) _2761_ : pout_data_stage0_0;
  assign _2763_ = rd_pout_data_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6997" *) data_hmult_stage0_in0 : pout_data_stage0_0;
  assign _1081_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6996" *) _2763_ : _2762_;
  assign _2764_ = rd_pout_data_stage0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6339" *) pout_mem_data_3 : pout_data_0_3;
  assign _2765_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6327" *) { data_8bit_7, data_8bit_6 } : { data_16bit_3[21], data_16bit_3[21], data_16bit_3[21], data_16bit_3[21], data_16bit_3[21], data_16bit_3[21], data_16bit_3 };
  assign _2766_ = rd_pout_data_stage0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6326" *) _2765_ : pout_data_0_3;
  assign _1080_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6325" *) _2766_ : _2764_;
  assign _2767_ = rd_pout_data_stage0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6339" *) pout_mem_data_2 : pout_data_0_2;
  assign _2768_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6327" *) { data_8bit_5, data_8bit_4 } : { data_16bit_2[21], data_16bit_2[21], data_16bit_2[21], data_16bit_2[21], data_16bit_2[21], data_16bit_2[21], data_16bit_2 };
  assign _2769_ = rd_pout_data_stage0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6326" *) _2768_ : pout_data_0_2;
  assign _1079_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6325" *) _2769_ : _2767_;
  assign _2770_ = rd_pout_data_stage0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6339" *) pout_mem_data_1 : pout_data_0_1;
  assign _2771_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6327" *) { data_8bit_3, data_8bit_2 } : { data_16bit_1[21], data_16bit_1[21], data_16bit_1[21], data_16bit_1[21], data_16bit_1[21], data_16bit_1[21], data_16bit_1 };
  assign _2772_ = rd_pout_data_stage0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6326" *) _2771_ : pout_data_0_1;
  assign _1078_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6325" *) _2772_ : _2770_;
  assign _2773_ = rd_pout_data_stage0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6339" *) pout_mem_data_0 : pout_data_0_0;
  assign _2774_ = int8_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6327" *) { data_8bit_1, data_8bit_0 } : { data_16bit_0[21], data_16bit_0[21], data_16bit_0[21], data_16bit_0[21], data_16bit_0[21], data_16bit_0[21], data_16bit_0 };
  assign _2775_ = rd_pout_data_stage0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6326" *) _2774_ : pout_data_0_0;
  assign _1077_ = _1828_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6325" *) _2775_ : _2773_;
  function [18:0] _5956_;
    input [18:0] a;
    input [132:0] b;
    input [6:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6284|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6277" *)
    (* parallel_case *)
    casez (s)
      7'b??????1:
        _5956_ = b[18:0];
      7'b?????1?:
        _5956_ = b[37:19];
      7'b????1??:
        _5956_ = b[56:38];
      7'b???1???:
        _5956_ = b[75:57];
      7'b??1????:
        _5956_ = b[94:76];
      7'b?1?????:
        _5956_ = b[113:95];
      7'b1??????:
        _5956_ = b[132:114];
      default:
        _5956_ = a;
    endcase
  endfunction
  assign pad_table_out = _5956_(19'b0000000000000000000, { reg2dp_pad_value_1x_cfg, reg2dp_pad_value_2x_cfg, reg2dp_pad_value_3x_cfg, reg2dp_pad_value_4x_cfg, reg2dp_pad_value_5x_cfg, reg2dp_pad_value_6x_cfg, reg2dp_pad_value_7x_cfg }, { _2782_, _2781_, _2780_, _2779_, _2778_, _2777_, _2776_ });
  assign _2776_ = pad_table_index == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6284|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6277" *) 3'b111;
  assign _2777_ = pad_table_index == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6283|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6277" *) 3'b110;
  assign _2778_ = pad_table_index == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6282|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6277" *) 3'b101;
  assign _2779_ = pad_table_index == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6281|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6277" *) 3'b100;
  assign _2780_ = pad_table_index == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6280|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6277" *) 2'b11;
  assign _2781_ = pad_table_index == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6279|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6277" *) 2'b10;
  assign _2782_ = pad_table_index == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6278|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6277" *) 1'b1;
  assign _1096_ = rd_pout_data_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6206" *) pout_mem_data[114:112] : pout_mem_size_v;
  assign _1095_ = rd_pout_data_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6206" *) pout_mem_data[111:84] : pout_mem_data_3;
  assign _1094_ = rd_pout_data_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6206" *) pout_mem_data[83:56] : pout_mem_data_2;
  assign _1093_ = rd_pout_data_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6206" *) pout_mem_data[55:28] : pout_mem_data_1;
  assign _1092_ = rd_pout_data_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6206" *) pout_mem_data[27:0] : pout_mem_data_0;
  function [114:0] _5969_;
    input [114:0] a;
    input [919:0] b;
    input [7:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6188|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6180" *)
    (* parallel_case *)
    casez (s)
      8'b???????1:
        _5969_ = b[114:0];
      8'b??????1?:
        _5969_ = b[229:115];
      8'b?????1??:
        _5969_ = b[344:230];
      8'b????1???:
        _5969_ = b[459:345];
      8'b???1????:
        _5969_ = b[574:460];
      8'b??1?????:
        _5969_ = b[689:575];
      8'b?1??????:
        _5969_ = b[804:690];
      8'b1???????:
        _5969_ = b[919:805];
      default:
        _5969_ = a;
    endcase
  endfunction
  assign pout_mem_data_act = _5969_(115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, { mem_data0[114:112], pooling_2d_result_0, mem_data1[114:112], pooling_2d_result_1, mem_data2[114:112], pooling_2d_result_2, mem_data3[114:112], pooling_2d_result_3, mem_data4[114:112], pooling_2d_result_4, mem_data5[114:112], pooling_2d_result_5, mem_data6[114:112], pooling_2d_result_6, mem_data7[114:112], pooling_2d_result_7 }, { _2790_, _2789_, _2788_, _2787_, _2786_, _2785_, _2784_, _2783_ });
  assign _2783_ = pout_mem_data_sel == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6188|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6180" *) 8'b10000000;
  assign _2784_ = pout_mem_data_sel == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6187|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6180" *) 7'b1000000;
  assign _2785_ = pout_mem_data_sel == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6186|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6180" *) 6'b100000;
  assign _2786_ = pout_mem_data_sel == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6185|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6180" *) 5'b10000;
  assign _2787_ = pout_mem_data_sel == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6184|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6180" *) 4'b1000;
  assign _2788_ = pout_mem_data_sel == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6183|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6180" *) 3'b100;
  assign _2789_ = pout_mem_data_sel == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6182|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6180" *) 2'b10;
  assign _2790_ = pout_mem_data_sel == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6181|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6180" *) 1'b1;
  assign _2791_ = pout_data_stage3_prdy ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6126" *) 1'b0 : pout_data_stage3_vld;
  assign _1091_ = pout_data_stage2_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6124" *) 1'b1 : _2791_;
  assign _1102_ = rd_pout_data_stage2_all ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6063" *) rd_pout_data_en_3d : rd_pout_data_en_4d;
  assign _1101_ = rd_pout_data_stage1_all ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6000" *) rd_pout_data_en_2d : rd_pout_data_en_3d;
  assign _2792_ = pout_data_stage2_prdy ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5991" *) 1'b0 : pout_data_stage2_vld;
  assign _1090_ = pout_data_stage1_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5989" *) 1'b1 : _2792_;
  assign _1100_ = load_wr_stage3_all ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5926" *) rd_pout_data_en_d : rd_pout_data_en_2d;
  assign _2793_ = pout_data_stage1_prdy ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5917" *) 1'b0 : pout_data_stage1_vld;
  assign _1089_ = wr_data_stage2_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5915" *) 1'b1 : _2793_;
  assign _1103_ = load_wr_stage2_all ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5852" *) rd_pout_data_en : rd_pout_data_en_d;
  assign _2794_ = _1773_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5837" *) _1264_[2:0] : rd_comb_lbuf_cnt;
  assign _1098_ = _2691_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5835" *) 3'b000 : _2794_;
  assign _2795_ = rd_sub_lbuf_end ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5824" *) _1263_ : rd_sub_lbuf_cnt;
  assign _1104_ = rd_comb_lbuf_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5822" *) 3'b000 : _2795_;
  assign _2796_ = rd_line_out ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5812" *) _1262_ : rd_line_out_cnt;
  assign _1099_ = _2690_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5810" *) 6'b000000 : _2796_;
  assign _1068_ = load_wr_stage2_all ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5706" *) one_width_disable_2d : one_width_disable_3d;
  assign _1013_ = load_wr_stage2_all ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5645" *) cur_datin_disable_2d : cur_datin_disable_3d;
  assign _1067_ = load_wr_stage1_all ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5584" *) one_width_disable_d : one_width_disable_2d;
  assign _1012_ = load_wr_stage1_all ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5523" *) cur_datin_disable_d : cur_datin_disable_2d;
  assign _1113_ = _2264_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5456" *) unit2d_cnt_pooling_last_d : unit2d_cnt_pooling_last_2d;
  assign _1062_ = _2263_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5395" *) mem_re_last_d : mem_re_last_2d;
  assign _1069_ = load_din_all ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5334" *) one_width_disable : one_width_disable_d;
  assign _1014_ = load_din_all ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5273" *) cur_datin_disable : cur_datin_disable_d;
  assign _1114_ = _2261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5212" *) unit2d_cnt_pooling_last : unit2d_cnt_pooling_last_d;
  assign _1063_ = _2262_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5151" *) mem_re_last : mem_re_last_d;
  assign _1017_ = _2261_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5090" *) flush_read_en : flush_read_en_d;
  assign _2797_ = unit2d_cnt_pooling_last_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5042" *) 3'b000 : _1261_;
  assign _2798_ = _1712_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5041" *) _2797_ : unit2d_cnt_pooling_last;
  assign _1112_ = wr_surface_dat_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5035" *) _2828_ : _2798_;
  assign _1057_ = wr_surface_dat_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5035" *) mem_re4_sel : mem_re4_sel_last;
  assign _1055_ = wr_surface_dat_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5035" *) mem_re3_sel : mem_re3_sel_last;
  assign _1053_ = wr_surface_dat_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5035" *) mem_re2_sel : mem_re2_sel_last;
  assign _1018_ = load_wr_stage2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4499" *) mem_raddr_2d : int_mem_waddr;
  assign _1027_ = load_wr_stage2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4438" *) mem_re_2d : int_mem_we;
  assign _1026_ = load_wr_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4421" *) { wr_line_end_2d, mem_data7[114:112], pooling_2d_result_7 } : int_mem_wdata_7;
  assign _1025_ = load_wr_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4421" *) { wr_line_end_2d, mem_data6[114:112], pooling_2d_result_6 } : int_mem_wdata_6;
  assign _1024_ = load_wr_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4421" *) { wr_line_end_2d, mem_data5[114:112], pooling_2d_result_5 } : int_mem_wdata_5;
  assign _1023_ = load_wr_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4421" *) { wr_line_end_2d, mem_data4[114:112], pooling_2d_result_4 } : int_mem_wdata_4;
  assign _1022_ = load_wr_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4421" *) { wr_line_end_2d, mem_data3[114:112], pooling_2d_result_3 } : int_mem_wdata_3;
  assign _1021_ = load_wr_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4421" *) { wr_line_end_2d, mem_data2[114:112], pooling_2d_result_2 } : int_mem_wdata_2;
  assign _1020_ = load_wr_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4421" *) { wr_line_end_2d, mem_data1[114:112], pooling_2d_result_1 } : int_mem_wdata_1;
  assign _1019_ = load_wr_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4421" *) { wr_line_end_2d, mem_data0[114:112], pooling_2d_result_0 } : int_mem_wdata_0;
  assign _2799_ = pout_data_stage0_prdy ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4372" *) 1'b0 : wr_data_stage2_vld;
  assign _1155_ = _1707_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4370" *) 1'b1 : _2799_;
  assign _2800_ = wr_data_stage1_prdy ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4358" *) 1'b0 : wr_data_stage1_vld;
  assign _1154_ = wr_data_stage0_vld ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4356" *) 1'b1 : _2800_;
  assign _2801_ = wr_data_stage0_prdy ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4343" *) 1'b0 : wr_data_stage0_vld;
  assign _1153_ = pooling1d_vld_rebuild ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4341" *) 1'b1 : _2801_;
  assign _1060_ = load_wr_stage1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4272" *) mem_re_d : mem_re_2d;
  assign _1061_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4211" *) mem_re : mem_re_d;
  assign _1050_ = _2252_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4148" *) sub_lbuf_dout_cnt : mem_raddr_d;
  assign _1058_ = load_wr_stage1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4087" *) mem_re_1st_d : mem_re_1st_2d;
  assign _1059_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4026" *) mem_re_1st : mem_re_1st_d;
  assign _1028_ = load_wr_stage1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3965" *) last_active_line_d : last_active_line_2d;
  assign _1029_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3904" *) active_last_line : last_active_line_d;
  assign _1162_ = load_wr_stage1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3843" *) wr_surface_dat_done_buf : wr_surface_dat_done_2d;
  assign _1049_ = load_wr_stage1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3782" *) mem_raddr_d : mem_raddr_2d;
  assign _1157_ = load_wr_stage1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3721" *) wr_line_end_buf : wr_line_end_2d;
  assign _1016_ = load_wr_stage1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3660" *) datin_buf : datin_buf_2d;
  assign _1047_ = load_wr_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3644" *) { unit2d_vsize_cnt_7_d, _3500_[111:0] } : mem_data7;
  assign _1045_ = load_wr_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3644" *) { unit2d_vsize_cnt_6_d, _3499_[111:0] } : mem_data6;
  assign _1043_ = load_wr_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3644" *) { unit2d_vsize_cnt_5_d, _3498_[111:0] } : mem_data5;
  assign _1041_ = load_wr_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3644" *) { unit2d_vsize_cnt_4_d, _3497_[111:0] } : mem_data4;
  assign _1039_ = load_wr_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3644" *) { unit2d_vsize_cnt_3_d, _3496_[111:0] } : mem_data3;
  assign _1037_ = load_wr_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3644" *) { unit2d_vsize_cnt_2_d, _3495_[111:0] } : mem_data2;
  assign _1035_ = load_wr_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3644" *) { unit2d_vsize_cnt_1_d, _3494_[111:0] } : mem_data1;
  assign _1033_ = load_wr_stage1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3644" *) { unit2d_vsize_cnt_0_d, _3493_[111:0] } : mem_data0;
  assign _1048_ = _1703_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3621" *) mem_rdata_7[114:0] : mem_data7_lst;
  assign _1046_ = _1703_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3621" *) mem_rdata_6[114:0] : mem_data6_lst;
  assign _1044_ = _1703_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3621" *) mem_rdata_5[114:0] : mem_data5_lst;
  assign _1042_ = _1703_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3621" *) mem_rdata_4[114:0] : mem_data4_lst;
  assign _1040_ = _1703_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3621" *) mem_rdata_3[114:0] : mem_data3_lst;
  assign _1038_ = _1703_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3621" *) mem_rdata_2[114:0] : mem_data2_lst;
  assign _1036_ = _1703_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3621" *) mem_rdata_1[114:0] : mem_data1_lst;
  assign _1034_ = _1703_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3621" *) mem_rdata_0[114:0] : mem_data0_lst;
  assign _2802_ = _2262_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3435" *) _1260_ : sub_lbuf_dout_cnt;
  assign _1107_ = _2637_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3432" *) 6'b000000 : _2802_;
  assign _2803_ = sub_lbuf_dout_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3422" *) _1259_ : wr_sub_lbuf_cnt;
  assign _1160_ = _2635_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3420" *) 3'b000 : _2803_;
  assign _1147_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3203" *) unit2d_vsize_7 : unit2d_vsize_cnt_7_d;
  assign _1145_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3142" *) unit2d_vsize_6 : unit2d_vsize_cnt_6_d;
  assign _1143_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3081" *) unit2d_vsize_5 : unit2d_vsize_cnt_5_d;
  assign _1141_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3020" *) unit2d_vsize_4 : unit2d_vsize_cnt_4_d;
  assign _1139_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2959" *) unit2d_vsize_3 : unit2d_vsize_cnt_3_d;
  assign _1137_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2898" *) unit2d_vsize_2 : unit2d_vsize_cnt_2_d;
  assign _1135_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2837" *) unit2d_vsize_1 : unit2d_vsize_cnt_1_d;
  assign _1133_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2776" *) unit2d_vsize_0 : unit2d_vsize_cnt_0_d;
  assign _2804_ = _1337_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2724" *) _1258_ : unit2d_vsize_cnt_7;
  assign _1146_ = unit2d_set[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2722" *) 3'b000 : _2804_;
  assign _2805_ = _1336_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2714" *) _1257_ : unit2d_vsize_cnt_6;
  assign _1144_ = unit2d_set[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2712" *) 3'b000 : _2805_;
  assign _2806_ = _1335_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2704" *) _1256_ : unit2d_vsize_cnt_5;
  assign _1142_ = unit2d_set[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2702" *) 3'b000 : _2806_;
  assign _2807_ = _1334_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2694" *) _1255_ : unit2d_vsize_cnt_4;
  assign _1140_ = unit2d_set[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2692" *) 3'b000 : _2807_;
  assign _2808_ = _1333_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2684" *) _1254_ : unit2d_vsize_cnt_3;
  assign _1138_ = unit2d_set[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2682" *) 3'b000 : _2808_;
  assign _2809_ = _1332_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2674" *) _1253_ : unit2d_vsize_cnt_2;
  assign _1136_ = unit2d_set[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2672" *) 3'b000 : _2809_;
  assign _2810_ = _1331_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2664" *) _1252_ : unit2d_vsize_cnt_1;
  assign _1134_ = unit2d_set[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2662" *) 3'b000 : _2810_;
  assign _2811_ = _1330_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2654" *) _1251_ : unit2d_vsize_cnt_0;
  assign _1132_ = unit2d_set[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2652" *) 3'b000 : _2811_;
  assign _1163_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2588" *) wr_surface_dat_done : wr_surface_dat_done_buf;
  assign _1158_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2527" *) wr_line_dat_done : wr_line_end_buf;
  assign _1015_ = load_din ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2466" *) pooling1d_pd : datin_buf;
  assign _2812_ = unit2d_clr[7] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2455" *) 1'b0 : unit2d_en[7];
  assign _2813_ = unit2d_set[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2453" *) 1'b1 : _2812_;
  assign _1123_ = wr_total_cube_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2451" *) 1'b0 : _2813_;
  assign _2814_ = unit2d_clr[6] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2439" *) 1'b0 : unit2d_en[6];
  assign _2815_ = unit2d_set[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2437" *) 1'b1 : _2814_;
  assign _1122_ = wr_total_cube_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2435" *) 1'b0 : _2815_;
  assign _2816_ = unit2d_clr[5] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2423" *) 1'b0 : unit2d_en[5];
  assign _2817_ = unit2d_set[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2421" *) 1'b1 : _2816_;
  assign _1121_ = wr_total_cube_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2419" *) 1'b0 : _2817_;
  assign _2818_ = unit2d_clr[4] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2407" *) 1'b0 : unit2d_en[4];
  assign _2819_ = unit2d_set[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2405" *) 1'b1 : _2818_;
  assign _1120_ = wr_total_cube_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2403" *) 1'b0 : _2819_;
  assign _2820_ = unit2d_clr[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2391" *) 1'b0 : unit2d_en[3];
  assign _2821_ = unit2d_set[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2389" *) 1'b1 : _2820_;
  assign _1119_ = wr_total_cube_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2387" *) 1'b0 : _2821_;
  assign _2822_ = unit2d_clr[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2375" *) 1'b0 : unit2d_en[2];
  assign _2823_ = unit2d_set[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2373" *) 1'b1 : _2822_;
  assign _1118_ = wr_total_cube_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2371" *) 1'b0 : _2823_;
  assign _2824_ = unit2d_clr[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2359" *) 1'b0 : unit2d_en[1];
  assign _2825_ = unit2d_set[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2357" *) 1'b1 : _2824_;
  assign _1117_ = wr_total_cube_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2355" *) 1'b0 : _2825_;
  assign _2826_ = unit2d_clr[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2343" *) 1'b0 : unit2d_en[0];
  assign _2827_ = unit2d_set[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2341" *) 1'b1 : _2826_;
  assign _1116_ = wr_total_cube_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2339" *) 1'b0 : _2827_;
  assign _2828_ = unit2d_cnt_pooling_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2314" *) 3'b000 : _1239_;
  assign _2829_ = _2623_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2313" *) _2828_ : unit2d_cnt_pooling;
  assign _1111_ = init_cnt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2311" *) 3'b000 : _2829_;
  assign _2830_ = stride_trig_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2299" *) 3'b000 : _1250_;
  assign _2831_ = stride_end ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2298" *) _2830_ : unit2d_cnt_stride;
  assign _1115_ = init_cnt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2296" *) padding_stride_num : _2831_;
  assign _2832_ = pooling1d_norm_rdy ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2279" *) _1249_ : one_width_bubble_cnt;
  assign _2833_ = one_width_bubble_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2277" *) 3'b000 : _2832_;
  assign _1065_ = one_width_disable ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2276" *) _2833_ : 3'b000;
  assign _2834_ = one_width_bubble_end ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2267" *) 1'b0 : one_width_disable;
  assign _1066_ = _1306_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2265" *) 1'b1 : _2834_;
  assign _1190_ = last_splitw ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2255" *) _2221_ : _3147_;
  assign _1166_ = first_splitw ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2253" *) _2220_ : _1190_;
  assign is_one_width_in = splitw_enable ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2251" *) _1166_ : _2219_;
  assign _2835_ = _2622_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2182" *) 3'b000 : _1248_;
  assign _2836_ = wr_line_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2181" *) _2835_ : last_out_cnt;
  assign _1030_ = last_out_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2180" *) _2836_ : 3'b000;
  assign _2837_ = last_out_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2169" *) 1'b0 : last_out_en;
  assign _2838_ = _2621_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2167" *) 1'b1 : _2837_;
  assign _1031_ = _2341_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2166" *) _2838_ : 1'b0;
  assign _2839_ = load_din ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2157" *) 1'b0 : cube_end_flag;
  assign _1010_ = wr_subcube_dat_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2155" *) 1'b1 : _2839_;
  assign _2840_ = line_end ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2139" *) _1247_ : bubble_cnt;
  assign _2841_ = bubble_en_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2137" *) 3'b000 : _2840_;
  assign _1004_ = cur_datin_disable ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2136" *) _2841_ : 3'b000;
  assign _2842_ = last_c ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2125" *) _1246_ : line_cnt;
  assign _2843_ = line_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2123" *) 13'b0000000000000 : _2842_;
  assign _1032_ = cur_datin_disable ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2122" *) _2843_ : 13'b0000000000000;
  assign _2844_ = one_width_norm_rdy ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2110" *) _1245_ : channel_cnt;
  assign _2845_ = last_c ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2107" *) 2'b00 : _2844_;
  assign _1009_ = cur_datin_disable ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2106" *) _2845_ : 2'b00;
  assign _1097_ = _2331_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2098" *) pout_width_cur : pout_width_cur_latch;
  assign _2846_ = bubble_en_end ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2080" *) 1'b0 : cur_datin_disable;
  assign _2847_ = _2620_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2078" *) 1'b1 : _2846_;
  assign _1011_ = _2619_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2076" *) 1'b1 : _2847_;
  assign _2848_ = one_width_bubble_end ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2067" *) 1'b0 : surfend_need_bubble_flg;
  assign _1110_ = _1292_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2065" *) 1'b1 : _2848_;
  assign _2849_ = one_width_bubble_end ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2057" *) 1'b0 : subend_need_flush_flg;
  assign _1108_ = _1290_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2055" *) 1'b1 : _2849_;
  assign _2850_ = _2205_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2021" *) 3'b101 : 3'b000;
  assign _2851_ = _2212_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2020" *) _2850_ : up_pnum5;
  assign _2852_ = _2210_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1994" *) 3'b000 : _2851_;
  assign _2853_ = _2208_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1974" *) 3'b000 : _2852_;
  assign _2854_ = _2206_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1954" *) 3'b000 : _2853_;
  assign _2855_ = _2204_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1940" *) 3'b000 : _2854_;
  assign _1152_ = _2203_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1934" *) 3'b000 : _2855_;
  assign _2856_ = _2205_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2021" *) 3'b100 : 3'b000;
  assign _2857_ = _2212_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2020" *) _2856_ : up_pnum4;
  assign _2858_ = _2210_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1994" *) _2856_ : _2857_;
  assign _2859_ = _2208_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1974" *) 3'b000 : _2858_;
  assign _2860_ = _2206_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1954" *) 3'b000 : _2859_;
  assign _2861_ = _2204_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1940" *) 3'b000 : _2860_;
  assign _1151_ = _2203_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1934" *) 3'b000 : _2861_;
  assign _2862_ = _2205_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2021" *) 2'b11 : 2'b00;
  assign _2863_ = _2212_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2020" *) _2862_ : up_pnum3;
  assign _2864_ = _2210_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1994" *) _2862_ : _2863_;
  assign _2865_ = _2208_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1974" *) _2862_ : _2864_;
  assign _2866_ = _2206_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1954" *) 2'b00 : _2865_;
  assign _2867_ = _2204_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1940" *) 2'b00 : _2866_;
  assign _1150_ = _2203_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1934" *) 2'b00 : _2867_;
  assign _2868_ = _2207_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2027" *) 2'b10 : 2'b00;
  assign _2869_ = _2205_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2021" *) 2'b10 : _2868_;
  assign _2870_ = _2212_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2020" *) _2869_ : up_pnum2;
  assign _2871_ = _2210_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1994" *) _2869_ : _2870_;
  assign _2872_ = _2205_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1975" *) 2'b10 : 2'b00;
  assign _2873_ = _2208_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1974" *) _2872_ : _2871_;
  assign _2874_ = _2206_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1954" *) _2872_ : _2873_;
  assign _2875_ = _2204_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1940" *) 2'b00 : _2874_;
  assign _1149_ = _2203_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1934" *) 2'b00 : _2875_;
  assign _2876_ = _2207_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2027" *) 1'b1 : _2618_;
  assign _2877_ = _2205_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2021" *) 1'b1 : _2876_;
  assign _2878_ = _2212_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2020" *) _2877_ : up_pnum1;
  assign _2879_ = _2207_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2001" *) 1'b1 : _2617_;
  assign _2880_ = _2205_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1995" *) 1'b1 : _2879_;
  assign _2881_ = _2210_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1994" *) _2880_ : _2878_;
  assign _2882_ = _2205_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1975" *) 1'b1 : _2616_;
  assign _2883_ = _2208_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1974" *) _2882_ : _2881_;
  assign _2884_ = _2205_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1955" *) 1'b1 : _2207_;
  assign _2885_ = _2206_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1954" *) _2884_ : _2883_;
  assign _2886_ = _2204_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1940" *) _2205_ : _2885_;
  assign _1148_ = _2203_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1934" *) 1'b0 : _2886_;
  assign _2887_ = _2202_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1918" *) unit2d_cnt_pooling_max : pnum_flush6;
  assign _2888_ = _2201_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1910" *) 3'b000 : _2887_;
  assign _2889_ = _2200_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1902" *) 3'b001 : _2888_;
  assign _2890_ = _2199_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1894" *) 3'b010 : _2889_;
  assign _2891_ = _2198_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1886" *) 3'b011 : _2890_;
  assign _2892_ = _2197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1878" *) 3'b100 : _2891_;
  assign _2893_ = _2196_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1870" *) 3'b101 : _2892_;
  assign _2894_ = unit2d_cnt_pooling_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1862" *) 3'b110 : _2893_;
  assign _1076_ = last_line_in ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1861" *) _2894_ : pnum_flush6;
  assign _2895_ = _2202_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1918" *) _1244_ : pnum_flush5;
  assign _2896_ = _2201_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1910" *) unit2d_cnt_pooling_max : _2895_;
  assign _2897_ = _2200_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1902" *) 3'b000 : _2896_;
  assign _2898_ = _2199_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1894" *) 3'b001 : _2897_;
  assign _2899_ = _2198_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1886" *) 3'b010 : _2898_;
  assign _2900_ = _2197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1878" *) 3'b011 : _2899_;
  assign _2901_ = _2196_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1870" *) 3'b100 : _2900_;
  assign _2902_ = unit2d_cnt_pooling_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1862" *) 3'b101 : _2901_;
  assign _1075_ = last_line_in ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1861" *) _2902_ : pnum_flush5;
  assign _2903_ = _2202_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1918" *) _1243_ : pnum_flush4;
  assign _2904_ = _2201_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1910" *) _1243_ : _2903_;
  assign _2905_ = _2200_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1902" *) unit2d_cnt_pooling_max : _2904_;
  assign _2906_ = _2199_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1894" *) 3'b000 : _2905_;
  assign _2907_ = _2198_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1886" *) 3'b001 : _2906_;
  assign _2908_ = _2197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1878" *) 3'b010 : _2907_;
  assign _2909_ = _2196_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1870" *) 3'b011 : _2908_;
  assign _2910_ = unit2d_cnt_pooling_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1862" *) 3'b100 : _2909_;
  assign _1074_ = last_line_in ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1861" *) _2910_ : pnum_flush4;
  assign _2911_ = _2202_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1918" *) _1242_ : pnum_flush3;
  assign _2912_ = _2201_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1910" *) _1242_ : _2911_;
  assign _2913_ = _2200_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1902" *) _1242_ : _2912_;
  assign _2914_ = _2199_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1894" *) unit2d_cnt_pooling_max : _2913_;
  assign _2915_ = _2198_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1886" *) 3'b000 : _2914_;
  assign _2916_ = _2197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1878" *) 3'b001 : _2915_;
  assign _2917_ = _2196_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1870" *) 3'b010 : _2916_;
  assign _2918_ = unit2d_cnt_pooling_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1862" *) 3'b011 : _2917_;
  assign _1073_ = last_line_in ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1861" *) _2918_ : pnum_flush3;
  assign _2919_ = _2202_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1918" *) _1241_ : pnum_flush2;
  assign _2920_ = _2201_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1910" *) _1241_ : _2919_;
  assign _2921_ = _2200_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1902" *) _1241_ : _2920_;
  assign _2922_ = _2199_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1894" *) _1241_ : _2921_;
  assign _2923_ = _2198_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1886" *) unit2d_cnt_pooling_max : _2922_;
  assign _2924_ = _2197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1878" *) 3'b000 : _2923_;
  assign _2925_ = _2196_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1870" *) 3'b001 : _2924_;
  assign _2926_ = unit2d_cnt_pooling_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1862" *) 3'b010 : _2925_;
  assign _1072_ = last_line_in ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1861" *) _2926_ : pnum_flush2;
  assign _2927_ = _2202_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1918" *) _1240_ : pnum_flush1;
  assign _2928_ = _2201_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1910" *) _1240_ : _2927_;
  assign _2929_ = _2200_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1902" *) _1240_ : _2928_;
  assign _2930_ = _2199_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1894" *) _1240_ : _2929_;
  assign _2931_ = _2198_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1886" *) _1240_ : _2930_;
  assign _2932_ = _2197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1878" *) unit2d_cnt_pooling_max : _2931_;
  assign _2933_ = _2196_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1870" *) 3'b000 : _2932_;
  assign _2934_ = unit2d_cnt_pooling_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1862" *) 3'b001 : _2933_;
  assign _1071_ = last_line_in ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1861" *) _2934_ : pnum_flush1;
  assign _2935_ = _2202_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1918" *) _1239_ : pnum_flush0;
  assign _2936_ = _2201_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1910" *) _1239_ : _2935_;
  assign _2937_ = _2200_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1902" *) _1239_ : _2936_;
  assign _2938_ = _2199_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1894" *) _1239_ : _2937_;
  assign _2939_ = _2198_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1886" *) _1239_ : _2938_;
  assign _2940_ = _2197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1878" *) _1239_ : _2939_;
  assign _2941_ = _2196_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1870" *) unit2d_cnt_pooling_max : _2940_;
  assign _2942_ = unit2d_cnt_pooling_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1862" *) 3'b000 : _2941_;
  assign _1070_ = last_line_in ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1861" *) _2942_ : pnum_flush0;
  assign _1915_[1:0] = _2611_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1839" *) 2'b10 : { 1'b0, _1914_[0] };
  assign _1916_[1:0] = _2606_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1837" *) 2'b11 : _1915_[1:0];
  assign _2943_ = _2601_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1835" *) 3'b100 : { 1'b0, _1916_[1:0] };
  assign _2944_ = _2596_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1833" *) 3'b101 : _2943_;
  assign _2945_ = _2591_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1831" *) 3'b110 : _2944_;
  assign _2946_ = _2586_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1829" *) 3'b111 : _2945_;
  assign _2947_ = _2033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1828" *) _2946_ : 3'b000;
  assign _1918_[1:0] = _2577_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1822" *) 2'b10 : { 1'b0, _1917_[0] };
  assign _1919_[1:0] = _2572_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1820" *) 2'b11 : _1918_[1:0];
  assign _2948_ = _2567_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1818" *) 3'b100 : { 1'b0, _1919_[1:0] };
  assign _2949_ = _2562_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1816" *) 3'b101 : _2948_;
  assign _2950_ = _2557_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1814" *) 3'b110 : _2949_;
  assign _2951_ = _2032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1813" *) _2950_ : _2947_;
  assign _1921_[1:0] = _2548_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1807" *) 2'b10 : { 1'b0, _1920_[0] };
  assign _1922_[1:0] = _2543_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1805" *) 2'b11 : _1921_[1:0];
  assign _2952_ = _2538_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1803" *) 3'b100 : { 1'b0, _1922_[1:0] };
  assign _2953_ = _2533_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1801" *) 3'b101 : _2952_;
  assign _2954_ = _2031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1800" *) _2953_ : _2951_;
  assign _1924_[1:0] = _2524_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1794" *) 2'b10 : { 1'b0, _1923_[0] };
  assign _1925_[1:0] = _2519_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1792" *) 2'b11 : _1924_[1:0];
  assign _2955_ = _2514_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1790" *) 3'b100 : { 1'b0, _1925_[1:0] };
  assign _2956_ = _2030_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1789" *) _2955_ : _2954_;
  assign _1927_[1:0] = _2505_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1783" *) 2'b10 : { 1'b0, _1926_[0] };
  assign _1928_[1:0] = _2500_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1781" *) 2'b11 : _1927_[1:0];
  assign _2957_ = _2029_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1780" *) { 1'b0, _1928_[1:0] } : _2956_;
  assign _1930_[1:0] = _2491_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1774" *) 2'b10 : { 1'b0, _1929_[0] };
  assign _1003_ = _2023_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1773" *) { 1'b0, _1930_[1:0] } : _2957_;
  assign next7_0 = _2033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1751" *) pnum_flush0 : 3'b000;
  assign next7_1 = _2033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1751" *) pnum_flush1 : 3'b000;
  assign next7_2 = _2033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1751" *) pnum_flush2 : 3'b000;
  assign next7_3 = _2033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1751" *) pnum_flush3 : 3'b000;
  assign next7_4 = _2033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1751" *) pnum_flush4 : 3'b000;
  assign next7_5 = _2033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1751" *) pnum_flush5 : 3'b000;
  assign next7_6 = _2033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1751" *) pnum_flush6 : 3'b000;
  assign _1181_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1717" *) pnum_flush0 : pnum_flush1;
  assign _1182_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1717" *) pnum_flush1 : pnum_flush2;
  assign _1183_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1717" *) pnum_flush2 : pnum_flush3;
  assign _1184_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1717" *) pnum_flush3 : pnum_flush4;
  assign _1185_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1717" *) pnum_flush4 : pnum_flush5;
  assign _1186_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1717" *) pnum_flush5 : pnum_flush6;
  assign next6_5 = _2032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1716" *) _1186_ : 3'b000;
  assign next6_4 = _2032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1716" *) _1185_ : 3'b000;
  assign next6_3 = _2032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1716" *) _1184_ : 3'b000;
  assign next6_2 = _2032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1716" *) _1183_ : 3'b000;
  assign next6_1 = _2032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1716" *) _1182_ : 3'b000;
  assign next6_0 = _2032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1716" *) _1181_ : 3'b000;
  assign _1200_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1684" *) pnum_flush1 : pnum_flush2;
  assign _1201_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1684" *) pnum_flush2 : pnum_flush3;
  assign _1202_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1684" *) pnum_flush3 : pnum_flush4;
  assign _1203_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1684" *) pnum_flush4 : pnum_flush5;
  assign _1204_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1684" *) pnum_flush5 : pnum_flush6;
  assign _1176_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1678" *) pnum_flush0 : _1200_;
  assign _1177_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1678" *) pnum_flush1 : _1201_;
  assign _1178_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1678" *) pnum_flush2 : _1202_;
  assign _1179_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1678" *) pnum_flush3 : _1203_;
  assign _1180_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1678" *) pnum_flush4 : _1204_;
  assign next5_4 = _2031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1677" *) _1180_ : 3'b000;
  assign next5_3 = _2031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1677" *) _1179_ : 3'b000;
  assign next5_2 = _2031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1677" *) _1178_ : 3'b000;
  assign next5_1 = _2031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1677" *) _1177_ : 3'b000;
  assign next5_0 = _2031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1677" *) _1176_ : 3'b000;
  assign _1213_ = _2026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1648" *) pnum_flush2 : pnum_flush3;
  assign _1214_ = _2026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1648" *) pnum_flush3 : pnum_flush4;
  assign _1215_ = _2026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1648" *) pnum_flush4 : pnum_flush5;
  assign _1216_ = _2026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1648" *) pnum_flush5 : pnum_flush6;
  assign _1196_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1643" *) pnum_flush1 : _1213_;
  assign _1197_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1643" *) pnum_flush2 : _1214_;
  assign _1198_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1643" *) pnum_flush3 : _1215_;
  assign _1199_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1643" *) pnum_flush4 : _1216_;
  assign _1172_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1638" *) pnum_flush0 : _1196_;
  assign _1173_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1638" *) pnum_flush1 : _1197_;
  assign _1174_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1638" *) pnum_flush2 : _1198_;
  assign _1175_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1638" *) pnum_flush3 : _1199_;
  assign next4_3 = _2030_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1637" *) _1175_ : 3'b000;
  assign next4_2 = _2030_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1637" *) _1174_ : 3'b000;
  assign next4_1 = _2030_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1637" *) _1173_ : 3'b000;
  assign next4_0 = _2030_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1637" *) _1172_ : 3'b000;
  assign _1221_ = _2027_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1611" *) pnum_flush3 : pnum_flush4;
  assign _1222_ = _2027_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1611" *) pnum_flush4 : pnum_flush5;
  assign _1223_ = _2027_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1611" *) pnum_flush5 : pnum_flush6;
  assign _1210_ = _2026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1607" *) pnum_flush2 : _1221_;
  assign _1211_ = _2026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1607" *) pnum_flush3 : _1222_;
  assign _1212_ = _2026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1607" *) pnum_flush4 : _1223_;
  assign _1193_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1603" *) pnum_flush1 : _1210_;
  assign _1194_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1603" *) pnum_flush2 : _1211_;
  assign _1195_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1603" *) pnum_flush3 : _1212_;
  assign _1169_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1599" *) pnum_flush0 : _1193_;
  assign _1170_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1599" *) pnum_flush1 : _1194_;
  assign _1171_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1599" *) pnum_flush2 : _1195_;
  assign next3_2 = _2029_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1598" *) _1171_ : 3'b000;
  assign next3_1 = _2029_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1598" *) _1170_ : 3'b000;
  assign next3_0 = _2029_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1598" *) _1169_ : 3'b000;
  assign _1226_ = _2028_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1575" *) pnum_flush4 : pnum_flush5;
  assign _1227_ = _2028_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1575" *) pnum_flush5 : pnum_flush6;
  assign _1219_ = _2027_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1572" *) pnum_flush3 : _1226_;
  assign _1220_ = _2027_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1572" *) pnum_flush4 : _1227_;
  assign _1208_ = _2026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1569" *) pnum_flush2 : _1219_;
  assign _1209_ = _2026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1569" *) pnum_flush3 : _1220_;
  assign _1191_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1566" *) pnum_flush1 : _1208_;
  assign _1192_ = _2025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1566" *) pnum_flush2 : _1209_;
  assign _1167_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1563" *) pnum_flush0 : _1191_;
  assign _1168_ = _2024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1563" *) pnum_flush1 : _1192_;
  assign next2_1 = _2023_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1562" *) _1168_ : 3'b000;
  assign next2_0 = _2023_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1562" *) _1167_ : 3'b000;
  assign _2958_ = _2288_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1541" *) _1237_ : 3'b000;
  assign _1005_ = pdp_op_start ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1540" *) _2958_ : bubble_num;
  assign _2959_ = _2960_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1523" *) bubble_add : 3'b000;
  assign _2961_ = _2288_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1520" *) _1238_ : _2959_;
  assign _2962_ = last_line_in ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1519" *) _2961_ : bubble_num_use;
  assign _2963_ = need_flush ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1512" *) flush_num : 3'b000;
  assign _1006_ = wr_subcube_dat_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1511" *) _2963_ : _2962_;
  assign _2964_ = _2288_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1520" *) 1'b1 : _2960_;
  assign _2965_ = last_line_in ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1519" *) _2964_ : need_bubble;
  assign _1064_ = wr_subcube_dat_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1511" *) need_flush : _2965_;
  assign _1164_ = small_active ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1488" *) samllH_flush_num : flush_num_cal;
  assign flush_num = _2022_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1486" *) 3'b000 : _1164_;
  assign _1224_ = _2021_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1473" *) 2'b10 : { 1'b0, _1228_ };
  assign _1217_ = _2020_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1471" *) 2'b11 : _1224_;
  assign _1205_ = _2019_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1469" *) 3'b100 : { 1'b0, _1217_ };
  assign _1187_ = _2018_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1467" *) 3'b101 : _1205_;
  assign samllH_flush_num = _2017_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1465" *) 3'b110 : _1187_;
  assign pad_r_remain = small_active ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1450" *) _3140_ : 6'b000000;
  assign _1229_[0] = _2338_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1434" *) 1'b0 : 1'b1;
  assign _1225_ = _2337_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1432" *) 2'b01 : { 1'b1, _1229_[0] };
  assign _1218_ = _2336_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1430" *) 2'b00 : _1225_;
  assign _1207_ = _2335_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1428" *) 3'b011 : { 1'b1, _1218_ };
  assign _1189_ = _2334_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1426" *) 3'b010 : _1207_;
  assign _1165_ = _2333_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1424" *) 3'b001 : _1189_;
  assign flush_num_cal = _2332_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1422" *) 3'b000 : _1165_;
  assign _2966_ = _2330_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1396" *) strip_ycnt_stride_f[2:0] : 3'b000;
  assign _2967_ = wr_line_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1393" *) _1236_[2:0] : strip_ycnt_psize;
  assign _2968_ = pooling_2d_rdy ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1391" *) pooling_size_minus_sride : _2967_;
  assign _2969_ = _2287_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1390" *) _2968_ : _2966_;
  assign _1105_ = init_cnt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1388" *) padding_v_cfg : _2969_;
  assign _1106_ = _2016_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1325" *) strip_ycnt_stride_f : strip_ycnt_stride;
  assign _1206_ = wr_line_dat_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1316" *) _1235_ : strip_ycnt_stride;
  assign _1188_ = stride_end ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1314" *) 4'b0000 : _1206_;
  assign strip_ycnt_stride_f = init_cnt ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1312" *) { 1'b0, strip_ycnt_offset } : _1188_;
  function [2:0] _6391_;
    input [2:0] a;
    input [8:0] b;
    input [2:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1295|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1292" *)
    (* parallel_case *)
    casez (s)
      3'b??1:
        _6391_ = b[2:0];
      3'b?1?:
        _6391_ = b[5:3];
      3'b1??:
        _6391_ = b[8:6];
      default:
        _6391_ = a;
    endcase
  endfunction
  assign padding_stride_num = _6391_({ 2'b00, padding_stride4_num[0] }, { padding_v_cfg, 1'b0, padding_v_cfg[2:1], 1'b0, padding_stride3_num }, { _2972_, _2971_, _2970_ });
  assign _2970_ = pooling_stride_v_cfg == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1295|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1292" *) 2'b10;
  assign _2971_ = pooling_stride_v_cfg == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1294|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1292" *) 1'b1;
  assign _2972_ = ! (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1293|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1292" *) pooling_stride_v_cfg;
  function [3:0] _6395_;
    input [3:0] a;
    input [11:0] b;
    input [2:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1265|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1262" *)
    (* parallel_case *)
    casez (s)
      3'b??1:
        _6395_ = b[3:0];
      3'b?1?:
        _6395_ = b[7:4];
      3'b1??:
        _6395_ = b[11:8];
      default:
        _6395_ = a;
    endcase
  endfunction
  assign bank_merge_num = _6395_(4'b0001, 12'b100001000010, { _1051_, _1052_, _2973_ });
  assign _2973_ = | (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1265|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1262" *) { _2248_, _2249_ };
  function [3:0] _6397_;
    input [3:0] a;
    input [11:0] b;
    input [2:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1251|./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1248" *)
    (* parallel_case *)
    casez (s)
      3'b??1:
        _6397_ = b[3:0];
      3'b?1?:
        _6397_ = b[7:4];
      3'b1??:
        _6397_ = b[11:8];
      default:
        _6397_ = a;
    endcase
  endfunction
  assign _2974_ = _6397_(4'b0010, { buffer_lines_0, buffer_lines_1, 3'b001, buffer_lines_2 }, { _2972_, _2971_, _2970_ });
  assign _2975_ = pooling_stride_big ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1245" *) 4'b0001 : _2974_;
  assign _1007_ = pdp_op_start ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1244" *) _2975_ : buffer_lines_num;
  assign _2976_ = wr_subcube_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1209" *) _1234_ : wr_splitc_cnt;
  assign _1159_ = wr_total_cube_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1207" *) 8'b00000000 : _2976_;
  assign _2977_ = wr_surface_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1197" *) _1233_[10:0] : surface_cnt_rd;
  assign _1109_ = wr_subcube_dat_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1195" *) 11'b00000000000 : _2977_;
  assign _2978_ = wr_line_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1176" *) _1232_ : wr_surface_dat_cnt;
  assign _1161_ = wr_surface_dat_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1174" *) 13'b0000000000000 : _2978_;
  assign _2979_ = stripe_receive_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1164" *) _1231_ : wr_line_dat_cnt;
  assign _1156_ = wr_line_dat_done ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1162" *) 13'b0000000000000 : _2979_;
  assign _1008_ = load_din ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1152" *) _1230_ : c_cnt;
  assign _2980_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3586" *) { datin_buf_2d[10], datin_buf_2d[11], datin_buf_2d[12], datin_buf_2d[13], datin_buf_2d[14] };
  assign _2981_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data0[10], mem_data0[11], mem_data0[12], mem_data0[13], mem_data0[14] };
  assign _2982_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data1[10], mem_data1[11], mem_data1[12], mem_data1[13], mem_data1[14] };
  assign _2983_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data2[10], mem_data2[11], mem_data2[12], mem_data2[13], mem_data2[14] };
  assign _2984_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data3[10], mem_data3[11], mem_data3[12], mem_data3[13], mem_data3[14] };
  assign _2985_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data4[10], mem_data4[11], mem_data4[12], mem_data4[13], mem_data4[14] };
  assign _2986_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data5[10], mem_data5[11], mem_data5[12], mem_data5[13], mem_data5[14] };
  assign _2987_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data6[10], mem_data6[11], mem_data6[12], mem_data6[13], mem_data6[14] };
  assign _2988_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data7[10], mem_data7[11], mem_data7[12], mem_data7[13], mem_data7[14] };
  assign _2989_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3588" *) { datin_buf_2d[38], datin_buf_2d[39], datin_buf_2d[40], datin_buf_2d[41], datin_buf_2d[42] };
  assign _2990_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data0[38], mem_data0[39], mem_data0[40], mem_data0[41], mem_data0[42] };
  assign _2991_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data1[38], mem_data1[39], mem_data1[40], mem_data1[41], mem_data1[42] };
  assign _2992_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data2[38], mem_data2[39], mem_data2[40], mem_data2[41], mem_data2[42] };
  assign _2993_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data3[38], mem_data3[39], mem_data3[40], mem_data3[41], mem_data3[42] };
  assign _2994_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data4[38], mem_data4[39], mem_data4[40], mem_data4[41], mem_data4[42] };
  assign _2995_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data5[38], mem_data5[39], mem_data5[40], mem_data5[41], mem_data5[42] };
  assign _2996_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data6[38], mem_data6[39], mem_data6[40], mem_data6[41], mem_data6[42] };
  assign _2997_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data7[38], mem_data7[39], mem_data7[40], mem_data7[41], mem_data7[42] };
  assign _2998_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3590" *) { datin_buf_2d[66], datin_buf_2d[67], datin_buf_2d[68], datin_buf_2d[69], datin_buf_2d[70] };
  assign _2999_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data0[66], mem_data0[67], mem_data0[68], mem_data0[69], mem_data0[70] };
  assign _3000_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data1[66], mem_data1[67], mem_data1[68], mem_data1[69], mem_data1[70] };
  assign _3001_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data2[66], mem_data2[67], mem_data2[68], mem_data2[69], mem_data2[70] };
  assign _3002_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data3[66], mem_data3[67], mem_data3[68], mem_data3[69], mem_data3[70] };
  assign _3003_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data4[66], mem_data4[67], mem_data4[68], mem_data4[69], mem_data4[70] };
  assign _3004_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data5[66], mem_data5[67], mem_data5[68], mem_data5[69], mem_data5[70] };
  assign _3005_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data6[66], mem_data6[67], mem_data6[68], mem_data6[69], mem_data6[70] };
  assign _3006_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data7[66], mem_data7[67], mem_data7[68], mem_data7[69], mem_data7[70] };
  assign _3007_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3592" *) { datin_buf_2d[94], datin_buf_2d[95], datin_buf_2d[96], datin_buf_2d[97], datin_buf_2d[98] };
  assign _3008_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data0[94], mem_data0[95], mem_data0[96], mem_data0[97], mem_data0[98] };
  assign _3009_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data1[94], mem_data1[95], mem_data1[96], mem_data1[97], mem_data1[98] };
  assign _3010_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data2[94], mem_data2[95], mem_data2[96], mem_data2[97], mem_data2[98] };
  assign _3011_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data3[94], mem_data3[95], mem_data3[96], mem_data3[97], mem_data3[98] };
  assign _3012_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data4[94], mem_data4[95], mem_data4[96], mem_data4[97], mem_data4[98] };
  assign _3013_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data5[94], mem_data5[95], mem_data5[96], mem_data5[97], mem_data5[98] };
  assign _3014_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data6[94], mem_data6[95], mem_data6[96], mem_data6[97], mem_data6[98] };
  assign _3015_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data7[94], mem_data7[95], mem_data7[96], mem_data7[97], mem_data7[98] };
  assign _3016_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7781" *) { fp16_4add_in_prdy[0], fp16_4add_in_prdy[1], fp16_4add_in_prdy[2], fp16_4add_in_prdy[3], fp16_4add_in_prdy[4], fp16_4add_in_prdy[5], fp16_4add_in_prdy[6], fp16_4add_in_prdy[7] };
  assign _3017_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7784" *) { fp16_4add_in_prdy[1], fp16_4add_in_prdy[2], fp16_4add_in_prdy[3], fp16_4add_in_prdy[4], fp16_4add_in_prdy[5], fp16_4add_in_prdy[6], fp16_4add_in_prdy[7] };
  assign _3018_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7785" *) { fp16_4add_in_prdy[0], fp16_4add_in_prdy[2], fp16_4add_in_prdy[3], fp16_4add_in_prdy[4], fp16_4add_in_prdy[5], fp16_4add_in_prdy[6], fp16_4add_in_prdy[7] };
  assign _3019_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7786" *) { fp16_4add_in_prdy[0], fp16_4add_in_prdy[1], fp16_4add_in_prdy[3], fp16_4add_in_prdy[4], fp16_4add_in_prdy[5], fp16_4add_in_prdy[6], fp16_4add_in_prdy[7] };
  assign _3020_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7787" *) { fp16_4add_in_prdy[0], fp16_4add_in_prdy[1], fp16_4add_in_prdy[2], fp16_4add_in_prdy[4], fp16_4add_in_prdy[5], fp16_4add_in_prdy[6], fp16_4add_in_prdy[7] };
  assign _3021_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7788" *) { fp16_4add_in_prdy[0], fp16_4add_in_prdy[1], fp16_4add_in_prdy[2], fp16_4add_in_prdy[3], fp16_4add_in_prdy[5], fp16_4add_in_prdy[6], fp16_4add_in_prdy[7] };
  assign _3022_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7789" *) { fp16_4add_in_prdy[0], fp16_4add_in_prdy[1], fp16_4add_in_prdy[2], fp16_4add_in_prdy[3], fp16_4add_in_prdy[4], fp16_4add_in_prdy[6], fp16_4add_in_prdy[7] };
  assign _3023_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7790" *) { fp16_4add_in_prdy[0], fp16_4add_in_prdy[1], fp16_4add_in_prdy[2], fp16_4add_in_prdy[3], fp16_4add_in_prdy[4], fp16_4add_in_prdy[5], fp16_4add_in_prdy[7] };
  assign _3024_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7791" *) { fp16_4add_in_prdy[0], fp16_4add_in_prdy[1], fp16_4add_in_prdy[2], fp16_4add_in_prdy[3], fp16_4add_in_prdy[4], fp16_4add_in_prdy[5], fp16_4add_in_prdy[6] };
  assign _3025_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7952" *) { fp16_4add_out_pvld[0], fp16_4add_out_pvld[1], fp16_4add_out_pvld[2], fp16_4add_out_pvld[3], fp16_4add_out_pvld[4], fp16_4add_out_pvld[5], fp16_4add_out_pvld[6], fp16_4add_out_pvld[7] };
  assign _3026_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7953" *) { fp16_4add_out_pvld[1], fp16_4add_out_pvld[2], fp16_4add_out_pvld[3], fp16_4add_out_pvld[4], fp16_4add_out_pvld[5], fp16_4add_out_pvld[6], fp16_4add_out_pvld[7] };
  assign _3027_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7954" *) { fp16_4add_out_pvld[0], fp16_4add_out_pvld[2], fp16_4add_out_pvld[3], fp16_4add_out_pvld[4], fp16_4add_out_pvld[5], fp16_4add_out_pvld[6], fp16_4add_out_pvld[7] };
  assign _3028_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7955" *) { fp16_4add_out_pvld[0], fp16_4add_out_pvld[1], fp16_4add_out_pvld[3], fp16_4add_out_pvld[4], fp16_4add_out_pvld[5], fp16_4add_out_pvld[6], fp16_4add_out_pvld[7] };
  assign _3029_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7956" *) { fp16_4add_out_pvld[0], fp16_4add_out_pvld[1], fp16_4add_out_pvld[2], fp16_4add_out_pvld[4], fp16_4add_out_pvld[5], fp16_4add_out_pvld[6], fp16_4add_out_pvld[7] };
  assign _3030_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7957" *) { fp16_4add_out_pvld[0], fp16_4add_out_pvld[1], fp16_4add_out_pvld[2], fp16_4add_out_pvld[3], fp16_4add_out_pvld[5], fp16_4add_out_pvld[6], fp16_4add_out_pvld[7] };
  assign _3031_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7958" *) { fp16_4add_out_pvld[0], fp16_4add_out_pvld[1], fp16_4add_out_pvld[2], fp16_4add_out_pvld[3], fp16_4add_out_pvld[4], fp16_4add_out_pvld[6], fp16_4add_out_pvld[7] };
  assign _3032_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7959" *) { fp16_4add_out_pvld[0], fp16_4add_out_pvld[1], fp16_4add_out_pvld[2], fp16_4add_out_pvld[3], fp16_4add_out_pvld[4], fp16_4add_out_pvld[5], fp16_4add_out_pvld[7] };
  assign _3033_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7960" *) { fp16_4add_out_pvld[0], fp16_4add_out_pvld[1], fp16_4add_out_pvld[2], fp16_4add_out_pvld[3], fp16_4add_out_pvld[4], fp16_4add_out_pvld[5], fp16_4add_out_pvld[6] };
  assign _3034_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8787" *) { fp16_mul_pad_line_rdy[0], fp16_mul_pad_line_rdy[1] };
  assign fp_mulw_prdy = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8849" *) { fp16_add_pad_in_a_rdy[0], fp16_add_pad_in_a_rdy[1], fp16_add_pad_in_a_rdy[2], fp16_add_pad_in_a_rdy[3], fp16_add_pad_in_b_rdy[0], fp16_add_pad_in_b_rdy[1], fp16_add_pad_in_b_rdy[2], fp16_add_pad_in_b_rdy[3] };
  assign _3035_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8850" *) { fp16_add_pad_in_a_rdy[1], fp16_add_pad_in_a_rdy[2], fp16_add_pad_in_a_rdy[3], fp16_add_pad_in_b_rdy[0], fp16_add_pad_in_b_rdy[1], fp16_add_pad_in_b_rdy[2], fp16_add_pad_in_b_rdy[3] };
  assign _3036_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8851" *) { fp16_add_pad_in_a_rdy[0], fp16_add_pad_in_a_rdy[2], fp16_add_pad_in_a_rdy[3], fp16_add_pad_in_b_rdy[0], fp16_add_pad_in_b_rdy[1], fp16_add_pad_in_b_rdy[2], fp16_add_pad_in_b_rdy[3] };
  assign _3037_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8852" *) { fp16_add_pad_in_a_rdy[0], fp16_add_pad_in_a_rdy[1], fp16_add_pad_in_a_rdy[3], fp16_add_pad_in_b_rdy[0], fp16_add_pad_in_b_rdy[1], fp16_add_pad_in_b_rdy[2], fp16_add_pad_in_b_rdy[3] };
  assign _3038_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8853" *) { fp16_add_pad_in_a_rdy[0], fp16_add_pad_in_a_rdy[1], fp16_add_pad_in_a_rdy[2], fp16_add_pad_in_b_rdy[0], fp16_add_pad_in_b_rdy[1], fp16_add_pad_in_b_rdy[2], fp16_add_pad_in_b_rdy[3] };
  assign _3039_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8854" *) { fp16_add_pad_in_a_rdy[0], fp16_add_pad_in_a_rdy[1], fp16_add_pad_in_a_rdy[2], fp16_add_pad_in_a_rdy[3], fp16_add_pad_in_b_rdy[1], fp16_add_pad_in_b_rdy[2], fp16_add_pad_in_b_rdy[3] };
  assign _3040_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8855" *) { fp16_add_pad_in_a_rdy[0], fp16_add_pad_in_a_rdy[1], fp16_add_pad_in_a_rdy[2], fp16_add_pad_in_a_rdy[3], fp16_add_pad_in_b_rdy[0], fp16_add_pad_in_b_rdy[2], fp16_add_pad_in_b_rdy[3] };
  assign _3041_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8856" *) { fp16_add_pad_in_a_rdy[0], fp16_add_pad_in_a_rdy[1], fp16_add_pad_in_a_rdy[2], fp16_add_pad_in_a_rdy[3], fp16_add_pad_in_b_rdy[0], fp16_add_pad_in_b_rdy[1], fp16_add_pad_in_b_rdy[3] };
  assign _3042_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8857" *) { fp16_add_pad_in_a_rdy[0], fp16_add_pad_in_a_rdy[1], fp16_add_pad_in_a_rdy[2], fp16_add_pad_in_a_rdy[3], fp16_add_pad_in_b_rdy[0], fp16_add_pad_in_b_rdy[1], fp16_add_pad_in_b_rdy[2] };
  assign _3043_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8910" *) { fp16_add_pad_out_vld[1], fp16_add_pad_out_vld[2], fp16_add_pad_out_vld[3] };
  assign _3044_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8911" *) { fp16_add_pad_out_vld[0], fp16_add_pad_out_vld[2], fp16_add_pad_out_vld[3] };
  assign _3045_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8912" *) { fp16_add_pad_out_vld[0], fp16_add_pad_out_vld[1], fp16_add_pad_out_vld[3] };
  assign _3046_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8913" *) { fp16_add_pad_out_vld[0], fp16_add_pad_out_vld[1], fp16_add_pad_out_vld[2] };
  assign fp16_add_pad_out_pvld = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8914" *) { fp16_add_pad_out_vld[0], fp16_add_pad_out_vld[1], fp16_add_pad_out_vld[2], fp16_add_pad_out_vld[3] };
  assign _3047_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8922" *) { fp16_mulw_in_a_rdy[1], fp16_mulw_in_a_rdy[2], fp16_mulw_in_a_rdy[3], fp16_mulw_in_b_rdy[0], fp16_mulw_in_b_rdy[1], fp16_mulw_in_b_rdy[2], fp16_mulw_in_b_rdy[3] };
  assign _3048_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8923" *) { fp16_mulw_in_a_rdy[0], fp16_mulw_in_a_rdy[2], fp16_mulw_in_a_rdy[3], fp16_mulw_in_b_rdy[0], fp16_mulw_in_b_rdy[1], fp16_mulw_in_b_rdy[2], fp16_mulw_in_b_rdy[3] };
  assign _3049_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8924" *) { fp16_mulw_in_a_rdy[0], fp16_mulw_in_a_rdy[1], fp16_mulw_in_a_rdy[3], fp16_mulw_in_b_rdy[0], fp16_mulw_in_b_rdy[1], fp16_mulw_in_b_rdy[2], fp16_mulw_in_b_rdy[3] };
  assign _3050_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8925" *) { fp16_mulw_in_a_rdy[0], fp16_mulw_in_a_rdy[1], fp16_mulw_in_a_rdy[2], fp16_mulw_in_b_rdy[0], fp16_mulw_in_b_rdy[1], fp16_mulw_in_b_rdy[2], fp16_mulw_in_b_rdy[3] };
  assign _3051_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8926" *) { fp16_mulw_in_a_rdy[0], fp16_mulw_in_a_rdy[1], fp16_mulw_in_a_rdy[2], fp16_mulw_in_a_rdy[3], fp16_mulw_in_b_rdy[1], fp16_mulw_in_b_rdy[2], fp16_mulw_in_b_rdy[3] };
  assign _3052_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8927" *) { fp16_mulw_in_a_rdy[0], fp16_mulw_in_a_rdy[1], fp16_mulw_in_a_rdy[2], fp16_mulw_in_a_rdy[3], fp16_mulw_in_b_rdy[0], fp16_mulw_in_b_rdy[2], fp16_mulw_in_b_rdy[3] };
  assign _3053_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8928" *) { fp16_mulw_in_a_rdy[0], fp16_mulw_in_a_rdy[1], fp16_mulw_in_a_rdy[2], fp16_mulw_in_a_rdy[3], fp16_mulw_in_b_rdy[0], fp16_mulw_in_b_rdy[1], fp16_mulw_in_b_rdy[3] };
  assign _3054_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8929" *) { fp16_mulw_in_a_rdy[0], fp16_mulw_in_a_rdy[1], fp16_mulw_in_a_rdy[2], fp16_mulw_in_a_rdy[3], fp16_mulw_in_b_rdy[0], fp16_mulw_in_b_rdy[1], fp16_mulw_in_b_rdy[2] };
  assign fp16_mulw_rdy = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8930" *) { fp16_mulw_in_a_rdy[0], fp16_mulw_in_a_rdy[1], fp16_mulw_in_a_rdy[2], fp16_mulw_in_a_rdy[3], fp16_mulw_in_b_rdy[0], fp16_mulw_in_b_rdy[1], fp16_mulw_in_b_rdy[2], fp16_mulw_in_b_rdy[3] };
  assign _3055_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8983" *) { fp16_mulw_out_vld[1], fp16_mulw_out_vld[2], fp16_mulw_out_vld[3] };
  assign _3056_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8984" *) { fp16_mulw_out_vld[0], fp16_mulw_out_vld[2], fp16_mulw_out_vld[3] };
  assign _3057_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8985" *) { fp16_mulw_out_vld[0], fp16_mulw_out_vld[1], fp16_mulw_out_vld[3] };
  assign _3058_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8986" *) { fp16_mulw_out_vld[0], fp16_mulw_out_vld[1], fp16_mulw_out_vld[2] };
  assign fp16_mulv_in_vld = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8988" *) { fp16_mulw_out_vld[0], fp16_mulw_out_vld[1], fp16_mulw_out_vld[2], fp16_mulw_out_vld[3] };
  assign _3059_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8994" *) { fp16_mulv_in_a_rdy[1], fp16_mulv_in_a_rdy[2], fp16_mulv_in_a_rdy[3], fp16_mulv_in_b_rdy[0], fp16_mulv_in_b_rdy[1], fp16_mulv_in_b_rdy[2], fp16_mulv_in_b_rdy[3] };
  assign _3060_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8995" *) { fp16_mulv_in_a_rdy[0], fp16_mulv_in_a_rdy[2], fp16_mulv_in_a_rdy[3], fp16_mulv_in_b_rdy[0], fp16_mulv_in_b_rdy[1], fp16_mulv_in_b_rdy[2], fp16_mulv_in_b_rdy[3] };
  assign _3061_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8996" *) { fp16_mulv_in_a_rdy[0], fp16_mulv_in_a_rdy[1], fp16_mulv_in_a_rdy[3], fp16_mulv_in_b_rdy[0], fp16_mulv_in_b_rdy[1], fp16_mulv_in_b_rdy[2], fp16_mulv_in_b_rdy[3] };
  assign _3062_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8997" *) { fp16_mulv_in_a_rdy[0], fp16_mulv_in_a_rdy[1], fp16_mulv_in_a_rdy[2], fp16_mulv_in_b_rdy[0], fp16_mulv_in_b_rdy[1], fp16_mulv_in_b_rdy[2], fp16_mulv_in_b_rdy[3] };
  assign _3063_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8998" *) { fp16_mulv_in_a_rdy[0], fp16_mulv_in_a_rdy[1], fp16_mulv_in_a_rdy[2], fp16_mulv_in_a_rdy[3], fp16_mulv_in_b_rdy[1], fp16_mulv_in_b_rdy[2], fp16_mulv_in_b_rdy[3] };
  assign _3064_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8999" *) { fp16_mulv_in_a_rdy[0], fp16_mulv_in_a_rdy[1], fp16_mulv_in_a_rdy[2], fp16_mulv_in_a_rdy[3], fp16_mulv_in_b_rdy[0], fp16_mulv_in_b_rdy[2], fp16_mulv_in_b_rdy[3] };
  assign _3065_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9000" *) { fp16_mulv_in_a_rdy[0], fp16_mulv_in_a_rdy[1], fp16_mulv_in_a_rdy[2], fp16_mulv_in_a_rdy[3], fp16_mulv_in_b_rdy[0], fp16_mulv_in_b_rdy[1], fp16_mulv_in_b_rdy[3] };
  assign _3066_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9001" *) { fp16_mulv_in_a_rdy[0], fp16_mulv_in_a_rdy[1], fp16_mulv_in_a_rdy[2], fp16_mulv_in_a_rdy[3], fp16_mulv_in_b_rdy[0], fp16_mulv_in_b_rdy[1], fp16_mulv_in_b_rdy[2] };
  assign fp16_mulv_rdy = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9002" *) { fp16_mulv_in_a_rdy[0], fp16_mulv_in_a_rdy[1], fp16_mulv_in_a_rdy[2], fp16_mulv_in_a_rdy[3], fp16_mulv_in_b_rdy[0], fp16_mulv_in_b_rdy[1], fp16_mulv_in_b_rdy[2], fp16_mulv_in_b_rdy[3] };
  assign _3067_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9099" *) { fp17T16_out_vld[1], fp17T16_out_vld[2], fp17T16_out_vld[3] };
  assign _3068_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9100" *) { fp17T16_out_vld[0], fp17T16_out_vld[2], fp17T16_out_vld[3] };
  assign _3069_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9101" *) { fp17T16_out_vld[0], fp17T16_out_vld[1], fp17T16_out_vld[3] };
  assign _3070_ = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9102" *) { fp17T16_out_vld[0], fp17T16_out_vld[1], fp17T16_out_vld[2] };
  assign fp_dp2wdma_pvld = & (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9104" *) { fp17T16_out_vld[0], fp17T16_out_vld[1], fp17T16_out_vld[2], fp17T16_out_vld[3] };
  assign _3071_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1186" *) { cube_out_channel[0], cube_out_channel[1], cube_out_channel[2], cube_out_channel[3] };
  assign _3072_[0] = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1189" *) { cube_out_channel[0], cube_out_channel[1], cube_out_channel[2], cube_out_channel[3], cube_out_channel[4] };
  assign _3073_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1440" *) { reg2dp_cube_in_height[3], reg2dp_cube_in_height[4], reg2dp_cube_in_height[5], reg2dp_cube_in_height[6], reg2dp_cube_in_height[7], reg2dp_cube_in_height[8], reg2dp_cube_in_height[9], reg2dp_cube_in_height[10], reg2dp_cube_in_height[11], reg2dp_cube_in_height[12] };
  assign _2960_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1523" *) { bubble_add[0], bubble_add[1], bubble_add[2] };
  assign _3074_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3586" *) { datin_buf_2d[0], datin_buf_2d[1], datin_buf_2d[2], datin_buf_2d[3], datin_buf_2d[4], datin_buf_2d[5], datin_buf_2d[6], datin_buf_2d[7], datin_buf_2d[8], datin_buf_2d[9] };
  assign _3075_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data0[0], mem_data0[1], mem_data0[2], mem_data0[3], mem_data0[4], mem_data0[5], mem_data0[6], mem_data0[7], mem_data0[8], mem_data0[9] };
  assign _3076_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data1[0], mem_data1[1], mem_data1[2], mem_data1[3], mem_data1[4], mem_data1[5], mem_data1[6], mem_data1[7], mem_data1[8], mem_data1[9] };
  assign _3077_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data2[0], mem_data2[1], mem_data2[2], mem_data2[3], mem_data2[4], mem_data2[5], mem_data2[6], mem_data2[7], mem_data2[8], mem_data2[9] };
  assign _3078_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data3[0], mem_data3[1], mem_data3[2], mem_data3[3], mem_data3[4], mem_data3[5], mem_data3[6], mem_data3[7], mem_data3[8], mem_data3[9] };
  assign _3079_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data4[0], mem_data4[1], mem_data4[2], mem_data4[3], mem_data4[4], mem_data4[5], mem_data4[6], mem_data4[7], mem_data4[8], mem_data4[9] };
  assign _3080_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data5[0], mem_data5[1], mem_data5[2], mem_data5[3], mem_data5[4], mem_data5[5], mem_data5[6], mem_data5[7], mem_data5[8], mem_data5[9] };
  assign _3081_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data6[0], mem_data6[1], mem_data6[2], mem_data6[3], mem_data6[4], mem_data6[5], mem_data6[6], mem_data6[7], mem_data6[8], mem_data6[9] };
  assign _3082_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3587" *) { mem_data7[0], mem_data7[1], mem_data7[2], mem_data7[3], mem_data7[4], mem_data7[5], mem_data7[6], mem_data7[7], mem_data7[8], mem_data7[9] };
  assign _3083_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3588" *) { datin_buf_2d[28], datin_buf_2d[29], datin_buf_2d[30], datin_buf_2d[31], datin_buf_2d[32], datin_buf_2d[33], datin_buf_2d[34], datin_buf_2d[35], datin_buf_2d[36], datin_buf_2d[37] };
  assign _3084_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data0[28], mem_data0[29], mem_data0[30], mem_data0[31], mem_data0[32], mem_data0[33], mem_data0[34], mem_data0[35], mem_data0[36], mem_data0[37] };
  assign _3085_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data1[28], mem_data1[29], mem_data1[30], mem_data1[31], mem_data1[32], mem_data1[33], mem_data1[34], mem_data1[35], mem_data1[36], mem_data1[37] };
  assign _3086_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data2[28], mem_data2[29], mem_data2[30], mem_data2[31], mem_data2[32], mem_data2[33], mem_data2[34], mem_data2[35], mem_data2[36], mem_data2[37] };
  assign _3087_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data3[28], mem_data3[29], mem_data3[30], mem_data3[31], mem_data3[32], mem_data3[33], mem_data3[34], mem_data3[35], mem_data3[36], mem_data3[37] };
  assign _3088_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data4[28], mem_data4[29], mem_data4[30], mem_data4[31], mem_data4[32], mem_data4[33], mem_data4[34], mem_data4[35], mem_data4[36], mem_data4[37] };
  assign _3089_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data5[28], mem_data5[29], mem_data5[30], mem_data5[31], mem_data5[32], mem_data5[33], mem_data5[34], mem_data5[35], mem_data5[36], mem_data5[37] };
  assign _3090_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data6[28], mem_data6[29], mem_data6[30], mem_data6[31], mem_data6[32], mem_data6[33], mem_data6[34], mem_data6[35], mem_data6[36], mem_data6[37] };
  assign _3091_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3589" *) { mem_data7[28], mem_data7[29], mem_data7[30], mem_data7[31], mem_data7[32], mem_data7[33], mem_data7[34], mem_data7[35], mem_data7[36], mem_data7[37] };
  assign _3092_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3590" *) { datin_buf_2d[56], datin_buf_2d[57], datin_buf_2d[58], datin_buf_2d[59], datin_buf_2d[60], datin_buf_2d[61], datin_buf_2d[62], datin_buf_2d[63], datin_buf_2d[64], datin_buf_2d[65] };
  assign _3093_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data0[56], mem_data0[57], mem_data0[58], mem_data0[59], mem_data0[60], mem_data0[61], mem_data0[62], mem_data0[63], mem_data0[64], mem_data0[65] };
  assign _3094_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data1[56], mem_data1[57], mem_data1[58], mem_data1[59], mem_data1[60], mem_data1[61], mem_data1[62], mem_data1[63], mem_data1[64], mem_data1[65] };
  assign _3095_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data2[56], mem_data2[57], mem_data2[58], mem_data2[59], mem_data2[60], mem_data2[61], mem_data2[62], mem_data2[63], mem_data2[64], mem_data2[65] };
  assign _3096_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data3[56], mem_data3[57], mem_data3[58], mem_data3[59], mem_data3[60], mem_data3[61], mem_data3[62], mem_data3[63], mem_data3[64], mem_data3[65] };
  assign _3097_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data4[56], mem_data4[57], mem_data4[58], mem_data4[59], mem_data4[60], mem_data4[61], mem_data4[62], mem_data4[63], mem_data4[64], mem_data4[65] };
  assign _3098_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data5[56], mem_data5[57], mem_data5[58], mem_data5[59], mem_data5[60], mem_data5[61], mem_data5[62], mem_data5[63], mem_data5[64], mem_data5[65] };
  assign _3099_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data6[56], mem_data6[57], mem_data6[58], mem_data6[59], mem_data6[60], mem_data6[61], mem_data6[62], mem_data6[63], mem_data6[64], mem_data6[65] };
  assign _3100_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3591" *) { mem_data7[56], mem_data7[57], mem_data7[58], mem_data7[59], mem_data7[60], mem_data7[61], mem_data7[62], mem_data7[63], mem_data7[64], mem_data7[65] };
  assign _3101_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3592" *) { datin_buf_2d[84], datin_buf_2d[85], datin_buf_2d[86], datin_buf_2d[87], datin_buf_2d[88], datin_buf_2d[89], datin_buf_2d[90], datin_buf_2d[91], datin_buf_2d[92], datin_buf_2d[93] };
  assign _3102_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data0[84], mem_data0[85], mem_data0[86], mem_data0[87], mem_data0[88], mem_data0[89], mem_data0[90], mem_data0[91], mem_data0[92], mem_data0[93] };
  assign _3103_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data1[84], mem_data1[85], mem_data1[86], mem_data1[87], mem_data1[88], mem_data1[89], mem_data1[90], mem_data1[91], mem_data1[92], mem_data1[93] };
  assign _3104_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data2[84], mem_data2[85], mem_data2[86], mem_data2[87], mem_data2[88], mem_data2[89], mem_data2[90], mem_data2[91], mem_data2[92], mem_data2[93] };
  assign _3105_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data3[84], mem_data3[85], mem_data3[86], mem_data3[87], mem_data3[88], mem_data3[89], mem_data3[90], mem_data3[91], mem_data3[92], mem_data3[93] };
  assign _3106_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data4[84], mem_data4[85], mem_data4[86], mem_data4[87], mem_data4[88], mem_data4[89], mem_data4[90], mem_data4[91], mem_data4[92], mem_data4[93] };
  assign _3107_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data5[84], mem_data5[85], mem_data5[86], mem_data5[87], mem_data5[88], mem_data5[89], mem_data5[90], mem_data5[91], mem_data5[92], mem_data5[93] };
  assign _3108_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data6[84], mem_data6[85], mem_data6[86], mem_data6[87], mem_data6[88], mem_data6[89], mem_data6[90], mem_data6[91], mem_data6[92], mem_data6[93] };
  assign _3109_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3593" *) { mem_data7[84], mem_data7[85], mem_data7[86], mem_data7[87], mem_data7[88], mem_data7[89], mem_data7[90], mem_data7[91], mem_data7[92], mem_data7[93] };
  assign _3110_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4148" *) { mem_re[0], mem_re[1], mem_re[2], mem_re[3], mem_re[4], mem_re[5], mem_re[6], mem_re[7] };
  assign _3111_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5090" *) { mem_re_last[0], mem_re_last[1], mem_re_last[2], mem_re_last[3], mem_re_last[4], mem_re_last[5], mem_re_last[6], mem_re_last[7] };
  assign _3112_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5456" *) { mem_re_last_d[0], mem_re_last_d[1], mem_re_last_d[2], mem_re_last_d[3], mem_re_last_d[4], mem_re_last_d[5], mem_re_last_d[6], mem_re_last_d[7] };
  assign rd_line_out = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5844" *) { pout_mem_data_sel[0], pout_mem_data_sel[1], pout_mem_data_sel[2], pout_mem_data_sel[3], pout_mem_data_sel[4], pout_mem_data_sel[5], pout_mem_data_sel[6], pout_mem_data_sel[7] };
  assign _3113_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5845" *) { mem_re_last_2d[0], mem_re_last_2d[1], mem_re_last_2d[2], mem_re_last_2d[3], mem_re_last_2d[4], mem_re_last_2d[5], mem_re_last_2d[6], mem_re_last_2d[7] };
  assign _3114_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6374" *) { data_hmult_16bit_0_ext[0], data_hmult_16bit_0_ext[1], data_hmult_16bit_0_ext[2], data_hmult_16bit_0_ext[3], data_hmult_16bit_0_ext[4], data_hmult_16bit_0_ext[5], data_hmult_16bit_0_ext[6], data_hmult_16bit_0_ext[7], data_hmult_16bit_0_ext[8], data_hmult_16bit_0_ext[9], data_hmult_16bit_0_ext[10], data_hmult_16bit_0_ext[11], data_hmult_16bit_0_ext[12], data_hmult_16bit_0_ext[13], data_hmult_16bit_0_ext[14] };
  assign _3115_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6375" *) { data_hmult_16bit_1_ext[0], data_hmult_16bit_1_ext[1], data_hmult_16bit_1_ext[2], data_hmult_16bit_1_ext[3], data_hmult_16bit_1_ext[4], data_hmult_16bit_1_ext[5], data_hmult_16bit_1_ext[6], data_hmult_16bit_1_ext[7], data_hmult_16bit_1_ext[8], data_hmult_16bit_1_ext[9], data_hmult_16bit_1_ext[10], data_hmult_16bit_1_ext[11], data_hmult_16bit_1_ext[12], data_hmult_16bit_1_ext[13], data_hmult_16bit_1_ext[14] };
  assign _3116_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6376" *) { data_hmult_16bit_2_ext[0], data_hmult_16bit_2_ext[1], data_hmult_16bit_2_ext[2], data_hmult_16bit_2_ext[3], data_hmult_16bit_2_ext[4], data_hmult_16bit_2_ext[5], data_hmult_16bit_2_ext[6], data_hmult_16bit_2_ext[7], data_hmult_16bit_2_ext[8], data_hmult_16bit_2_ext[9], data_hmult_16bit_2_ext[10], data_hmult_16bit_2_ext[11], data_hmult_16bit_2_ext[12], data_hmult_16bit_2_ext[13], data_hmult_16bit_2_ext[14] };
  assign _3117_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6377" *) { data_hmult_16bit_3_ext[0], data_hmult_16bit_3_ext[1], data_hmult_16bit_3_ext[2], data_hmult_16bit_3_ext[3], data_hmult_16bit_3_ext[4], data_hmult_16bit_3_ext[5], data_hmult_16bit_3_ext[6], data_hmult_16bit_3_ext[7], data_hmult_16bit_3_ext[8], data_hmult_16bit_3_ext[9], data_hmult_16bit_3_ext[10], data_hmult_16bit_3_ext[11], data_hmult_16bit_3_ext[12], data_hmult_16bit_3_ext[13], data_hmult_16bit_3_ext[14] };
  assign _3118_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6587" *) { data_hmult_8bit_0_lsb_ext[0], data_hmult_8bit_0_lsb_ext[1], data_hmult_8bit_0_lsb_ext[2], data_hmult_8bit_0_lsb_ext[3], data_hmult_8bit_0_lsb_ext[4], data_hmult_8bit_0_lsb_ext[5], data_hmult_8bit_0_lsb_ext[6], data_hmult_8bit_0_lsb_ext[7], data_hmult_8bit_0_lsb_ext[8], data_hmult_8bit_0_lsb_ext[9], data_hmult_8bit_0_lsb_ext[10], data_hmult_8bit_0_lsb_ext[11], data_hmult_8bit_0_lsb_ext[12], data_hmult_8bit_0_lsb_ext[13], data_hmult_8bit_0_lsb_ext[14] };
  assign _3119_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6588" *) { data_hmult_8bit_0_msb_ext[0], data_hmult_8bit_0_msb_ext[1], data_hmult_8bit_0_msb_ext[2], data_hmult_8bit_0_msb_ext[3], data_hmult_8bit_0_msb_ext[4], data_hmult_8bit_0_msb_ext[5], data_hmult_8bit_0_msb_ext[6], data_hmult_8bit_0_msb_ext[7], data_hmult_8bit_0_msb_ext[8], data_hmult_8bit_0_msb_ext[9], data_hmult_8bit_0_msb_ext[10], data_hmult_8bit_0_msb_ext[11], data_hmult_8bit_0_msb_ext[12], data_hmult_8bit_0_msb_ext[13], data_hmult_8bit_0_msb_ext[14] };
  assign _3120_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6589" *) { data_hmult_8bit_1_lsb_ext[0], data_hmult_8bit_1_lsb_ext[1], data_hmult_8bit_1_lsb_ext[2], data_hmult_8bit_1_lsb_ext[3], data_hmult_8bit_1_lsb_ext[4], data_hmult_8bit_1_lsb_ext[5], data_hmult_8bit_1_lsb_ext[6], data_hmult_8bit_1_lsb_ext[7], data_hmult_8bit_1_lsb_ext[8], data_hmult_8bit_1_lsb_ext[9], data_hmult_8bit_1_lsb_ext[10], data_hmult_8bit_1_lsb_ext[11], data_hmult_8bit_1_lsb_ext[12], data_hmult_8bit_1_lsb_ext[13], data_hmult_8bit_1_lsb_ext[14] };
  assign _3121_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6590" *) { data_hmult_8bit_1_msb_ext[0], data_hmult_8bit_1_msb_ext[1], data_hmult_8bit_1_msb_ext[2], data_hmult_8bit_1_msb_ext[3], data_hmult_8bit_1_msb_ext[4], data_hmult_8bit_1_msb_ext[5], data_hmult_8bit_1_msb_ext[6], data_hmult_8bit_1_msb_ext[7], data_hmult_8bit_1_msb_ext[8], data_hmult_8bit_1_msb_ext[9], data_hmult_8bit_1_msb_ext[10], data_hmult_8bit_1_msb_ext[11], data_hmult_8bit_1_msb_ext[12], data_hmult_8bit_1_msb_ext[13], data_hmult_8bit_1_msb_ext[14] };
  assign _3122_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6591" *) { data_hmult_8bit_2_lsb_ext[0], data_hmult_8bit_2_lsb_ext[1], data_hmult_8bit_2_lsb_ext[2], data_hmult_8bit_2_lsb_ext[3], data_hmult_8bit_2_lsb_ext[4], data_hmult_8bit_2_lsb_ext[5], data_hmult_8bit_2_lsb_ext[6], data_hmult_8bit_2_lsb_ext[7], data_hmult_8bit_2_lsb_ext[8], data_hmult_8bit_2_lsb_ext[9], data_hmult_8bit_2_lsb_ext[10], data_hmult_8bit_2_lsb_ext[11], data_hmult_8bit_2_lsb_ext[12], data_hmult_8bit_2_lsb_ext[13], data_hmult_8bit_2_lsb_ext[14] };
  assign _3123_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6592" *) { data_hmult_8bit_2_msb_ext[0], data_hmult_8bit_2_msb_ext[1], data_hmult_8bit_2_msb_ext[2], data_hmult_8bit_2_msb_ext[3], data_hmult_8bit_2_msb_ext[4], data_hmult_8bit_2_msb_ext[5], data_hmult_8bit_2_msb_ext[6], data_hmult_8bit_2_msb_ext[7], data_hmult_8bit_2_msb_ext[8], data_hmult_8bit_2_msb_ext[9], data_hmult_8bit_2_msb_ext[10], data_hmult_8bit_2_msb_ext[11], data_hmult_8bit_2_msb_ext[12], data_hmult_8bit_2_msb_ext[13], data_hmult_8bit_2_msb_ext[14] };
  assign _3124_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6593" *) { data_hmult_8bit_3_lsb_ext[0], data_hmult_8bit_3_lsb_ext[1], data_hmult_8bit_3_lsb_ext[2], data_hmult_8bit_3_lsb_ext[3], data_hmult_8bit_3_lsb_ext[4], data_hmult_8bit_3_lsb_ext[5], data_hmult_8bit_3_lsb_ext[6], data_hmult_8bit_3_lsb_ext[7], data_hmult_8bit_3_lsb_ext[8], data_hmult_8bit_3_lsb_ext[9], data_hmult_8bit_3_lsb_ext[10], data_hmult_8bit_3_lsb_ext[11], data_hmult_8bit_3_lsb_ext[12], data_hmult_8bit_3_lsb_ext[13], data_hmult_8bit_3_lsb_ext[14] };
  assign _3125_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6594" *) { data_hmult_8bit_3_msb_ext[0], data_hmult_8bit_3_msb_ext[1], data_hmult_8bit_3_msb_ext[2], data_hmult_8bit_3_msb_ext[3], data_hmult_8bit_3_msb_ext[4], data_hmult_8bit_3_msb_ext[5], data_hmult_8bit_3_msb_ext[6], data_hmult_8bit_3_msb_ext[7], data_hmult_8bit_3_msb_ext[8], data_hmult_8bit_3_msb_ext[9], data_hmult_8bit_3_msb_ext[10], data_hmult_8bit_3_msb_ext[11], data_hmult_8bit_3_msb_ext[12], data_hmult_8bit_3_msb_ext[13], data_hmult_8bit_3_msb_ext[14] };
  assign _3126_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7029" *) { data_vmult_16bit_0_ext[0], data_vmult_16bit_0_ext[1], data_vmult_16bit_0_ext[2], data_vmult_16bit_0_ext[3], data_vmult_16bit_0_ext[4], data_vmult_16bit_0_ext[5], data_vmult_16bit_0_ext[6], data_vmult_16bit_0_ext[7], data_vmult_16bit_0_ext[8], data_vmult_16bit_0_ext[9], data_vmult_16bit_0_ext[10], data_vmult_16bit_0_ext[11], data_vmult_16bit_0_ext[12], data_vmult_16bit_0_ext[13], data_vmult_16bit_0_ext[14] };
  assign _3127_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7030" *) { data_vmult_16bit_1_ext[0], data_vmult_16bit_1_ext[1], data_vmult_16bit_1_ext[2], data_vmult_16bit_1_ext[3], data_vmult_16bit_1_ext[4], data_vmult_16bit_1_ext[5], data_vmult_16bit_1_ext[6], data_vmult_16bit_1_ext[7], data_vmult_16bit_1_ext[8], data_vmult_16bit_1_ext[9], data_vmult_16bit_1_ext[10], data_vmult_16bit_1_ext[11], data_vmult_16bit_1_ext[12], data_vmult_16bit_1_ext[13], data_vmult_16bit_1_ext[14] };
  assign _3128_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7031" *) { data_vmult_16bit_2_ext[0], data_vmult_16bit_2_ext[1], data_vmult_16bit_2_ext[2], data_vmult_16bit_2_ext[3], data_vmult_16bit_2_ext[4], data_vmult_16bit_2_ext[5], data_vmult_16bit_2_ext[6], data_vmult_16bit_2_ext[7], data_vmult_16bit_2_ext[8], data_vmult_16bit_2_ext[9], data_vmult_16bit_2_ext[10], data_vmult_16bit_2_ext[11], data_vmult_16bit_2_ext[12], data_vmult_16bit_2_ext[13], data_vmult_16bit_2_ext[14] };
  assign _3129_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7032" *) { data_vmult_16bit_3_ext[0], data_vmult_16bit_3_ext[1], data_vmult_16bit_3_ext[2], data_vmult_16bit_3_ext[3], data_vmult_16bit_3_ext[4], data_vmult_16bit_3_ext[5], data_vmult_16bit_3_ext[6], data_vmult_16bit_3_ext[7], data_vmult_16bit_3_ext[8], data_vmult_16bit_3_ext[9], data_vmult_16bit_3_ext[10], data_vmult_16bit_3_ext[11], data_vmult_16bit_3_ext[12], data_vmult_16bit_3_ext[13], data_vmult_16bit_3_ext[14] };
  assign _3130_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7242" *) { data_vmult_8bit_0_lsb_ext[0], data_vmult_8bit_0_lsb_ext[1], data_vmult_8bit_0_lsb_ext[2], data_vmult_8bit_0_lsb_ext[3], data_vmult_8bit_0_lsb_ext[4], data_vmult_8bit_0_lsb_ext[5], data_vmult_8bit_0_lsb_ext[6], data_vmult_8bit_0_lsb_ext[7], data_vmult_8bit_0_lsb_ext[8], data_vmult_8bit_0_lsb_ext[9], data_vmult_8bit_0_lsb_ext[10], data_vmult_8bit_0_lsb_ext[11], data_vmult_8bit_0_lsb_ext[12], data_vmult_8bit_0_lsb_ext[13], data_vmult_8bit_0_lsb_ext[14] };
  assign _3131_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7243" *) { data_vmult_8bit_0_msb_ext[0], data_vmult_8bit_0_msb_ext[1], data_vmult_8bit_0_msb_ext[2], data_vmult_8bit_0_msb_ext[3], data_vmult_8bit_0_msb_ext[4], data_vmult_8bit_0_msb_ext[5], data_vmult_8bit_0_msb_ext[6], data_vmult_8bit_0_msb_ext[7], data_vmult_8bit_0_msb_ext[8], data_vmult_8bit_0_msb_ext[9], data_vmult_8bit_0_msb_ext[10], data_vmult_8bit_0_msb_ext[11], data_vmult_8bit_0_msb_ext[12], data_vmult_8bit_0_msb_ext[13], data_vmult_8bit_0_msb_ext[14] };
  assign _3132_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7244" *) { data_vmult_8bit_1_lsb_ext[0], data_vmult_8bit_1_lsb_ext[1], data_vmult_8bit_1_lsb_ext[2], data_vmult_8bit_1_lsb_ext[3], data_vmult_8bit_1_lsb_ext[4], data_vmult_8bit_1_lsb_ext[5], data_vmult_8bit_1_lsb_ext[6], data_vmult_8bit_1_lsb_ext[7], data_vmult_8bit_1_lsb_ext[8], data_vmult_8bit_1_lsb_ext[9], data_vmult_8bit_1_lsb_ext[10], data_vmult_8bit_1_lsb_ext[11], data_vmult_8bit_1_lsb_ext[12], data_vmult_8bit_1_lsb_ext[13], data_vmult_8bit_1_lsb_ext[14] };
  assign _3133_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7245" *) { data_vmult_8bit_1_msb_ext[0], data_vmult_8bit_1_msb_ext[1], data_vmult_8bit_1_msb_ext[2], data_vmult_8bit_1_msb_ext[3], data_vmult_8bit_1_msb_ext[4], data_vmult_8bit_1_msb_ext[5], data_vmult_8bit_1_msb_ext[6], data_vmult_8bit_1_msb_ext[7], data_vmult_8bit_1_msb_ext[8], data_vmult_8bit_1_msb_ext[9], data_vmult_8bit_1_msb_ext[10], data_vmult_8bit_1_msb_ext[11], data_vmult_8bit_1_msb_ext[12], data_vmult_8bit_1_msb_ext[13], data_vmult_8bit_1_msb_ext[14] };
  assign _3134_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7246" *) { data_vmult_8bit_2_lsb_ext[0], data_vmult_8bit_2_lsb_ext[1], data_vmult_8bit_2_lsb_ext[2], data_vmult_8bit_2_lsb_ext[3], data_vmult_8bit_2_lsb_ext[4], data_vmult_8bit_2_lsb_ext[5], data_vmult_8bit_2_lsb_ext[6], data_vmult_8bit_2_lsb_ext[7], data_vmult_8bit_2_lsb_ext[8], data_vmult_8bit_2_lsb_ext[9], data_vmult_8bit_2_lsb_ext[10], data_vmult_8bit_2_lsb_ext[11], data_vmult_8bit_2_lsb_ext[12], data_vmult_8bit_2_lsb_ext[13], data_vmult_8bit_2_lsb_ext[14] };
  assign _3135_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7247" *) { data_vmult_8bit_2_msb_ext[0], data_vmult_8bit_2_msb_ext[1], data_vmult_8bit_2_msb_ext[2], data_vmult_8bit_2_msb_ext[3], data_vmult_8bit_2_msb_ext[4], data_vmult_8bit_2_msb_ext[5], data_vmult_8bit_2_msb_ext[6], data_vmult_8bit_2_msb_ext[7], data_vmult_8bit_2_msb_ext[8], data_vmult_8bit_2_msb_ext[9], data_vmult_8bit_2_msb_ext[10], data_vmult_8bit_2_msb_ext[11], data_vmult_8bit_2_msb_ext[12], data_vmult_8bit_2_msb_ext[13], data_vmult_8bit_2_msb_ext[14] };
  assign _3136_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7248" *) { data_vmult_8bit_3_lsb_ext[0], data_vmult_8bit_3_lsb_ext[1], data_vmult_8bit_3_lsb_ext[2], data_vmult_8bit_3_lsb_ext[3], data_vmult_8bit_3_lsb_ext[4], data_vmult_8bit_3_lsb_ext[5], data_vmult_8bit_3_lsb_ext[6], data_vmult_8bit_3_lsb_ext[7], data_vmult_8bit_3_lsb_ext[8], data_vmult_8bit_3_lsb_ext[9], data_vmult_8bit_3_lsb_ext[10], data_vmult_8bit_3_lsb_ext[11], data_vmult_8bit_3_lsb_ext[12], data_vmult_8bit_3_lsb_ext[13], data_vmult_8bit_3_lsb_ext[14] };
  assign _3137_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7249" *) { data_vmult_8bit_3_msb_ext[0], data_vmult_8bit_3_msb_ext[1], data_vmult_8bit_3_msb_ext[2], data_vmult_8bit_3_msb_ext[3], data_vmult_8bit_3_msb_ext[4], data_vmult_8bit_3_msb_ext[5], data_vmult_8bit_3_msb_ext[6], data_vmult_8bit_3_msb_ext[7], data_vmult_8bit_3_msb_ext[8], data_vmult_8bit_3_msb_ext[9], data_vmult_8bit_3_msb_ext[10], data_vmult_8bit_3_msb_ext[11], data_vmult_8bit_3_msb_ext[12], data_vmult_8bit_3_msb_ext[13], data_vmult_8bit_3_msb_ext[14] };
  assign _3138_ = | (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8762" *) { _2732_[0], _2732_[1], _2732_[2], _2732_[3], _2732_[4], _2732_[5], _2732_[6], _2732_[7] };
  assign { _3139_[31], _3139_[9:0] } = surface_num - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1201" *) 1'b1;
  assign strip_ycnt_offset = padding_v_cfg - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1299" *) _1913_[2:0];
  assign pooling_size_minus_sride = pooling_size_v_cfg - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1383" *) pooling_stride_v_cfg[2:0];
  assign _3140_ = h_pt_pb - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1451" *) reg2dp_kernel_height;
  assign _1931_[3:0] = buffer_lines_0 - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1504" *) padding_v_cfg;
  assign _3141_ = flush_num - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1522" *) first_out_num[2:0];
  assign flush_in_next_surf = flush_num - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1549" *) bubble_num;
  assign bubble_num_dec = bubble_num_use - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2146" *) 1'b1;
  assign _3142_ = flush_num - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2175" *) bubble_num_use;
  assign first_out_num_dec2 = _3142_ - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2175" *) 1'b1;
  assign flush_num_dec1 = flush_num - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2191" *) 1'b1;
  assign unit2d_cnt_pooling_max = buffer_lines_num[2:0] - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2322" *) 1'b1;
  assign rest_height = reg2dp_cube_in_height - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2326" *) wr_surface_dat_cnt;
  assign { _3143_[31], _3143_[3:0] } = bank_merge_num - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3426" *) 1'b1;
  assign { _3144_[31], _3144_[3:0] } = buffer_lines_num - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5841" *) 1'b1;
  assign pad_table_index = pooling_size_v_cfg - (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6221" *) pout_mem_size_v_use;
  assign surface_num = int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1190" *) surface_num_1 : surface_num_0;
  assign _3145_[9:0] = first_splitw ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1222" *) pooling_out_fwidth_cfg : pooling_out_mwidth_cfg;
  assign _3146_[9:0] = last_splitw ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1222" *) pooling_out_lwidth_cfg : _3145_[9:0];
  assign pout_width_cur = splitw_enable ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1222" *) { 3'b000, _3146_[9:0] } : reg2dp_cube_out_width;
  assign buffer_lines_2 = _2284_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1236" *) 1'b0 : 1'b1;
  assign padding_stride3_num = _2285_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1280" *) 2'b10 : { 1'b0, _2286_ };
  assign first_out_num = small_active ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:1504" *) cube_in_height_cfg : _1931_[3:0];
  assign _3147_ = _2297_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2258" *) _2222_ : 1'b0;
  assign unit2d_vsize1_0 = mem_re1_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2729" *) unit2d_vsize_cnt_0 : 3'b000;
  assign unit2d_vsize2_0 = mem_re2_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2738" *) unit2d_vsize_cnt_0 : 3'b000;
  assign unit2d_vsize2_4 = mem_re2_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2742" *) unit2d_vsize_cnt_1 : 3'b000;
  assign unit2d_vsize3_0 = mem_re3_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2747" *) unit2d_vsize_cnt_0 : 3'b000;
  assign unit2d_vsize3_2 = mem_re3_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2749" *) unit2d_vsize_cnt_1 : 3'b000;
  assign unit2d_vsize3_4 = mem_re3_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2751" *) unit2d_vsize_cnt_2 : 3'b000;
  assign unit2d_vsize3_6 = mem_re3_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2753" *) unit2d_vsize_cnt_3 : 3'b000;
  assign unit2d_vsize4_0 = mem_re4_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2756" *) unit2d_vsize_cnt_0 : 3'b000;
  assign unit2d_vsize4_1 = mem_re4_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2757" *) unit2d_vsize_cnt_1 : 3'b000;
  assign unit2d_vsize4_2 = mem_re4_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2758" *) unit2d_vsize_cnt_2 : 3'b000;
  assign unit2d_vsize4_3 = mem_re4_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2759" *) unit2d_vsize_cnt_3 : 3'b000;
  assign unit2d_vsize4_4 = mem_re4_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2760" *) unit2d_vsize_cnt_4 : 3'b000;
  assign unit2d_vsize4_5 = mem_re4_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2761" *) unit2d_vsize_cnt_5 : 3'b000;
  assign unit2d_vsize4_6 = mem_re4_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2762" *) unit2d_vsize_cnt_6 : 3'b000;
  assign unit2d_vsize4_7 = mem_re4_sel ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:2763" *) unit2d_vsize_cnt_7 : 3'b000;
  assign _3148_ = wr_line_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3274" *) 1'b0 : unit2d_mem_1strd[0];
  assign _1124_ = unit2d_set[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3274" *) 1'b1 : _3148_;
  assign _3149_ = wr_line_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3281" *) 1'b0 : unit2d_mem_1strd[1];
  assign _1125_ = unit2d_set[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3281" *) 1'b1 : _3149_;
  assign _3150_ = wr_line_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3288" *) 1'b0 : unit2d_mem_1strd[2];
  assign _1126_ = unit2d_set[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3288" *) 1'b1 : _3150_;
  assign _3151_ = wr_line_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3295" *) 1'b0 : unit2d_mem_1strd[3];
  assign _1127_ = unit2d_set[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3295" *) 1'b1 : _3151_;
  assign _3152_ = wr_line_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3302" *) 1'b0 : unit2d_mem_1strd[4];
  assign _1128_ = unit2d_set[4] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3302" *) 1'b1 : _3152_;
  assign _3153_ = wr_line_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3309" *) 1'b0 : unit2d_mem_1strd[5];
  assign _1129_ = unit2d_set[5] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3309" *) 1'b1 : _3153_;
  assign _3154_ = wr_line_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3316" *) 1'b0 : unit2d_mem_1strd[6];
  assign _1130_ = unit2d_set[6] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3316" *) 1'b1 : _3154_;
  assign _3155_ = wr_line_dat_done ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3323" *) 1'b0 : unit2d_mem_1strd[7];
  assign _1131_ = unit2d_set[7] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3323" *) 1'b1 : _3155_;
  assign { _0001_, _0000_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3472" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign { _0101_, _0100_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3472" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign { _0201_, _0200_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3472" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign { _0301_, _0300_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3472" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign { _0003_, _0002_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data0[27:0] : 28'b0000000000000000000000000000;
  assign { _0103_, _0102_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data0[55:28] : 28'b0000000000000000000000000000;
  assign { _0203_, _0202_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data0[83:56] : 28'b0000000000000000000000000000;
  assign { _0303_, _0302_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data0[111:84] : 28'b0000000000000000000000000000;
  assign { _0017_, _0016_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data1[27:0] : 28'b0000000000000000000000000000;
  assign { _0117_, _0116_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data1[55:28] : 28'b0000000000000000000000000000;
  assign { _0217_, _0216_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data1[83:56] : 28'b0000000000000000000000000000;
  assign { _0317_, _0316_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data1[111:84] : 28'b0000000000000000000000000000;
  assign { _0029_, _0028_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data2[27:0] : 28'b0000000000000000000000000000;
  assign { _0129_, _0128_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data2[55:28] : 28'b0000000000000000000000000000;
  assign { _0229_, _0228_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data2[83:56] : 28'b0000000000000000000000000000;
  assign { _0329_, _0328_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data2[111:84] : 28'b0000000000000000000000000000;
  assign { _0041_, _0040_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data3[27:0] : 28'b0000000000000000000000000000;
  assign { _0141_, _0140_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data3[55:28] : 28'b0000000000000000000000000000;
  assign { _0241_, _0240_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data3[83:56] : 28'b0000000000000000000000000000;
  assign { _0341_, _0340_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data3[111:84] : 28'b0000000000000000000000000000;
  assign { _0053_, _0052_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data4[27:0] : 28'b0000000000000000000000000000;
  assign { _0153_, _0152_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data4[55:28] : 28'b0000000000000000000000000000;
  assign { _0253_, _0252_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data4[83:56] : 28'b0000000000000000000000000000;
  assign { _0353_, _0352_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data4[111:84] : 28'b0000000000000000000000000000;
  assign { _0065_, _0064_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data5[27:0] : 28'b0000000000000000000000000000;
  assign { _0165_, _0164_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data5[55:28] : 28'b0000000000000000000000000000;
  assign { _0265_, _0264_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data5[83:56] : 28'b0000000000000000000000000000;
  assign { _0365_, _0364_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data5[111:84] : 28'b0000000000000000000000000000;
  assign { _0077_, _0076_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data6[27:0] : 28'b0000000000000000000000000000;
  assign { _0177_, _0176_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data6[55:28] : 28'b0000000000000000000000000000;
  assign { _0277_, _0276_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data6[83:56] : 28'b0000000000000000000000000000;
  assign { _0377_, _0376_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data6[111:84] : 28'b0000000000000000000000000000;
  assign { _0089_, _0088_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data7[27:0] : 28'b0000000000000000000000000000;
  assign { _0189_, _0188_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data7[55:28] : 28'b0000000000000000000000000000;
  assign { _0289_, _0288_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data7[83:56] : 28'b0000000000000000000000000000;
  assign { _0389_, _0388_ } = reg2dp_int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3473" *) mem_data7[111:84] : 28'b0000000000000000000000000000;
  assign _0006_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3474" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign _0106_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3474" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign _0206_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3474" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign _0306_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3474" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign _0007_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data0[27:0] : 28'b0000000000000000000000000000;
  assign _0107_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data0[55:28] : 28'b0000000000000000000000000000;
  assign _0207_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data0[83:56] : 28'b0000000000000000000000000000;
  assign _0307_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data0[111:84] : 28'b0000000000000000000000000000;
  assign _0019_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data1[27:0] : 28'b0000000000000000000000000000;
  assign _0119_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data1[55:28] : 28'b0000000000000000000000000000;
  assign _0219_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data1[83:56] : 28'b0000000000000000000000000000;
  assign _0319_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data1[111:84] : 28'b0000000000000000000000000000;
  assign _0031_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data2[27:0] : 28'b0000000000000000000000000000;
  assign _0131_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data2[55:28] : 28'b0000000000000000000000000000;
  assign _0231_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data2[83:56] : 28'b0000000000000000000000000000;
  assign _0331_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data2[111:84] : 28'b0000000000000000000000000000;
  assign _0043_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data3[27:0] : 28'b0000000000000000000000000000;
  assign _0143_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data3[55:28] : 28'b0000000000000000000000000000;
  assign _0243_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data3[83:56] : 28'b0000000000000000000000000000;
  assign _0343_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data3[111:84] : 28'b0000000000000000000000000000;
  assign _0055_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data4[27:0] : 28'b0000000000000000000000000000;
  assign _0155_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data4[55:28] : 28'b0000000000000000000000000000;
  assign _0255_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data4[83:56] : 28'b0000000000000000000000000000;
  assign _0355_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data4[111:84] : 28'b0000000000000000000000000000;
  assign _0067_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data5[27:0] : 28'b0000000000000000000000000000;
  assign _0167_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data5[55:28] : 28'b0000000000000000000000000000;
  assign _0267_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data5[83:56] : 28'b0000000000000000000000000000;
  assign _0367_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data5[111:84] : 28'b0000000000000000000000000000;
  assign _0079_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data6[27:0] : 28'b0000000000000000000000000000;
  assign _0179_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data6[55:28] : 28'b0000000000000000000000000000;
  assign _0279_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data6[83:56] : 28'b0000000000000000000000000000;
  assign _0379_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data6[111:84] : 28'b0000000000000000000000000000;
  assign _0091_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data7[27:0] : 28'b0000000000000000000000000000;
  assign _0191_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data7[55:28] : 28'b0000000000000000000000000000;
  assign _0291_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data7[83:56] : 28'b0000000000000000000000000000;
  assign _0391_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3475" *) mem_data7[111:84] : 28'b0000000000000000000000000000;
  assign _0004_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3476" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign _0104_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3476" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign _0204_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3476" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign _0304_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3476" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign _0005_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data0[27:0] : 28'b0000000000000000000000000000;
  assign _0105_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data0[55:28] : 28'b0000000000000000000000000000;
  assign _0205_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data0[83:56] : 28'b0000000000000000000000000000;
  assign _0305_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data0[111:84] : 28'b0000000000000000000000000000;
  assign _0018_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data1[27:0] : 28'b0000000000000000000000000000;
  assign _0118_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data1[55:28] : 28'b0000000000000000000000000000;
  assign _0218_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data1[83:56] : 28'b0000000000000000000000000000;
  assign _0318_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data1[111:84] : 28'b0000000000000000000000000000;
  assign _0030_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data2[27:0] : 28'b0000000000000000000000000000;
  assign _0130_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data2[55:28] : 28'b0000000000000000000000000000;
  assign _0230_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data2[83:56] : 28'b0000000000000000000000000000;
  assign _0330_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data2[111:84] : 28'b0000000000000000000000000000;
  assign _0042_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data3[27:0] : 28'b0000000000000000000000000000;
  assign _0142_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data3[55:28] : 28'b0000000000000000000000000000;
  assign _0242_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data3[83:56] : 28'b0000000000000000000000000000;
  assign _0342_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data3[111:84] : 28'b0000000000000000000000000000;
  assign _0054_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data4[27:0] : 28'b0000000000000000000000000000;
  assign _0154_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data4[55:28] : 28'b0000000000000000000000000000;
  assign _0254_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data4[83:56] : 28'b0000000000000000000000000000;
  assign _0354_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data4[111:84] : 28'b0000000000000000000000000000;
  assign _0066_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data5[27:0] : 28'b0000000000000000000000000000;
  assign _0166_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data5[55:28] : 28'b0000000000000000000000000000;
  assign _0266_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data5[83:56] : 28'b0000000000000000000000000000;
  assign _0366_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data5[111:84] : 28'b0000000000000000000000000000;
  assign _0078_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data6[27:0] : 28'b0000000000000000000000000000;
  assign _0178_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data6[55:28] : 28'b0000000000000000000000000000;
  assign _0278_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data6[83:56] : 28'b0000000000000000000000000000;
  assign _0378_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data6[111:84] : 28'b0000000000000000000000000000;
  assign _0090_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data7[27:0] : 28'b0000000000000000000000000000;
  assign _0190_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data7[55:28] : 28'b0000000000000000000000000000;
  assign _0290_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data7[83:56] : 28'b0000000000000000000000000000;
  assign _0390_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3477" *) mem_data7[111:84] : 28'b0000000000000000000000000000;
  assign _0402_ = _1367_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0000_ : _0002_;
  assign _0466_ = _1368_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0100_ : _0102_;
  assign _0530_ = _1369_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0200_ : _0202_;
  assign _0594_ = _1370_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0300_ : _0302_;
  assign _0410_ = _1371_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0000_ : _0016_;
  assign _0474_ = _1372_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0100_ : _0116_;
  assign _0538_ = _1373_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0200_ : _0216_;
  assign _0602_ = _1374_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0300_ : _0316_;
  assign _0418_ = _1375_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0000_ : _0028_;
  assign _0482_ = _1376_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0100_ : _0128_;
  assign _0546_ = _1377_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0200_ : _0228_;
  assign _0610_ = _1378_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0300_ : _0328_;
  assign _0426_ = _1379_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0000_ : _0040_;
  assign _0490_ = _1380_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0100_ : _0140_;
  assign _0554_ = _1381_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0200_ : _0240_;
  assign _0618_ = _1382_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0300_ : _0340_;
  assign _0434_ = _1383_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0000_ : _0052_;
  assign _0498_ = _1384_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0100_ : _0152_;
  assign _0562_ = _1385_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0200_ : _0252_;
  assign _0626_ = _1386_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0300_ : _0352_;
  assign _0442_ = _1387_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0000_ : _0064_;
  assign _0506_ = _1388_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0100_ : _0164_;
  assign _0570_ = _1389_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0200_ : _0264_;
  assign _0634_ = _1390_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0300_ : _0364_;
  assign _0450_ = _1391_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0000_ : _0076_;
  assign _0514_ = _1392_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0100_ : _0176_;
  assign _0578_ = _1393_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0200_ : _0276_;
  assign _0642_ = _1394_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0300_ : _0376_;
  assign _0458_ = _1395_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0000_ : _0088_;
  assign _0522_ = _1396_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0100_ : _0188_;
  assign _0586_ = _1397_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0200_ : _0288_;
  assign _0650_ = _1398_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3481" *) _0300_ : _0388_;
  assign _0404_ = _1399_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0001_ : _0003_;
  assign _0468_ = _1400_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0101_ : _0103_;
  assign _0532_ = _1401_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0201_ : _0203_;
  assign _0596_ = _1402_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0301_ : _0303_;
  assign _0412_ = _1403_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0001_ : _0017_;
  assign _0476_ = _1404_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0101_ : _0117_;
  assign _0540_ = _1405_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0201_ : _0217_;
  assign _0604_ = _1406_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0301_ : _0317_;
  assign _0420_ = _1407_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0001_ : _0029_;
  assign _0484_ = _1408_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0101_ : _0129_;
  assign _0548_ = _1409_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0201_ : _0229_;
  assign _0612_ = _1410_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0301_ : _0329_;
  assign _0428_ = _1411_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0001_ : _0041_;
  assign _0492_ = _1412_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0101_ : _0141_;
  assign _0556_ = _1413_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0201_ : _0241_;
  assign _0620_ = _1414_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0301_ : _0341_;
  assign _0436_ = _1415_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0001_ : _0053_;
  assign _0500_ = _1416_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0101_ : _0153_;
  assign _0564_ = _1417_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0201_ : _0253_;
  assign _0628_ = _1418_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0301_ : _0353_;
  assign _0444_ = _1419_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0001_ : _0065_;
  assign _0508_ = _1420_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0101_ : _0165_;
  assign _0572_ = _1421_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0201_ : _0265_;
  assign _0636_ = _1422_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0301_ : _0365_;
  assign _0452_ = _1423_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0001_ : _0077_;
  assign _0516_ = _1424_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0101_ : _0177_;
  assign _0580_ = _1425_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0201_ : _0277_;
  assign _0644_ = _1426_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0301_ : _0377_;
  assign _0460_ = _1427_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0001_ : _0089_;
  assign _0524_ = _1428_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0101_ : _0189_;
  assign _0588_ = _1429_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0201_ : _0289_;
  assign _0652_ = _1430_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3482" *) _0301_ : _0389_;
  assign _0400_ = _1431_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0006_ : _0007_;
  assign _0464_ = _1432_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0106_ : _0107_;
  assign _0528_ = _1433_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0206_ : _0207_;
  assign _0592_ = _1434_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0306_ : _0307_;
  assign _0408_ = _1435_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0006_ : _0019_;
  assign _0472_ = _1436_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0106_ : _0119_;
  assign _0536_ = _1437_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0206_ : _0219_;
  assign _0600_ = _1438_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0306_ : _0319_;
  assign _0416_ = _1439_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0006_ : _0031_;
  assign _0480_ = _1440_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0106_ : _0131_;
  assign _0544_ = _1441_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0206_ : _0231_;
  assign _0608_ = _1442_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0306_ : _0331_;
  assign _0424_ = _1443_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0006_ : _0043_;
  assign _0488_ = _1444_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0106_ : _0143_;
  assign _0552_ = _1445_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0206_ : _0243_;
  assign _0616_ = _1446_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0306_ : _0343_;
  assign _0432_ = _1447_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0006_ : _0055_;
  assign _0496_ = _1448_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0106_ : _0155_;
  assign _0560_ = _1449_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0206_ : _0255_;
  assign _0624_ = _1450_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0306_ : _0355_;
  assign _0440_ = _1451_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0006_ : _0067_;
  assign _0504_ = _1452_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0106_ : _0167_;
  assign _0568_ = _1453_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0206_ : _0267_;
  assign _0632_ = _1454_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0306_ : _0367_;
  assign _0448_ = _1455_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0006_ : _0079_;
  assign _0512_ = _1456_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0106_ : _0179_;
  assign _0576_ = _1457_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0206_ : _0279_;
  assign _0640_ = _1458_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0306_ : _0379_;
  assign _0456_ = _1459_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0006_ : _0091_;
  assign _0520_ = _1460_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0106_ : _0191_;
  assign _0584_ = _1461_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0206_ : _0291_;
  assign _0648_ = _1462_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3483" *) _0306_ : _0391_;
  assign _3156_ = _2298_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0005_ : _0004_;
  assign _3157_ = _2299_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0105_ : _0104_;
  assign _3158_ = _2300_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0205_ : _0204_;
  assign _3159_ = _2301_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0305_ : _0304_;
  assign _3160_ = _2302_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0018_ : _0004_;
  assign _3161_ = _2303_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0118_ : _0104_;
  assign _3162_ = _2304_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0218_ : _0204_;
  assign _3163_ = _2305_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0318_ : _0304_;
  assign _3164_ = _2306_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0030_ : _0004_;
  assign _3165_ = _2307_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0130_ : _0104_;
  assign _3166_ = _2308_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0230_ : _0204_;
  assign _3167_ = _2309_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0330_ : _0304_;
  assign _3168_ = _2310_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0042_ : _0004_;
  assign _3169_ = _2311_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0142_ : _0104_;
  assign _3170_ = _2312_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0242_ : _0204_;
  assign _3171_ = _2313_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0342_ : _0304_;
  assign _3172_ = _2314_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0054_ : _0004_;
  assign _3173_ = _2315_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0154_ : _0104_;
  assign _3174_ = _2316_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0254_ : _0204_;
  assign _3175_ = _2317_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0354_ : _0304_;
  assign _3176_ = _2318_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0066_ : _0004_;
  assign _3177_ = _2319_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0166_ : _0104_;
  assign _3178_ = _2320_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0266_ : _0204_;
  assign _3179_ = _2321_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0366_ : _0304_;
  assign _3180_ = _2322_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0078_ : _0004_;
  assign _3181_ = _2323_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0178_ : _0104_;
  assign _3182_ = _2324_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0278_ : _0204_;
  assign _3183_ = _2325_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0378_ : _0304_;
  assign _3184_ = _2326_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0090_ : _0004_;
  assign _3185_ = _2327_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0190_ : _0104_;
  assign _3186_ = _2328_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0290_ : _0204_;
  assign _3187_ = _2329_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3484" *) _0390_ : _0304_;
  assign _3188_ = _2298_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0004_ : _0005_;
  assign _3189_ = _2299_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0104_ : _0105_;
  assign _3190_ = _2300_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0204_ : _0205_;
  assign _3191_ = _2301_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0304_ : _0305_;
  assign _3192_ = _2302_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0004_ : _0018_;
  assign _3193_ = _2303_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0104_ : _0118_;
  assign _3194_ = _2304_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0204_ : _0218_;
  assign _3195_ = _2305_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0304_ : _0318_;
  assign _3196_ = _2306_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0004_ : _0030_;
  assign _3197_ = _2307_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0104_ : _0130_;
  assign _3198_ = _2308_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0204_ : _0230_;
  assign _3199_ = _2309_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0304_ : _0330_;
  assign _3200_ = _2310_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0004_ : _0042_;
  assign _3201_ = _2311_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0104_ : _0142_;
  assign _3202_ = _2312_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0204_ : _0242_;
  assign _3203_ = _2313_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0304_ : _0342_;
  assign _3204_ = _2314_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0004_ : _0054_;
  assign _3205_ = _2315_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0104_ : _0154_;
  assign _3206_ = _2316_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0204_ : _0254_;
  assign _3207_ = _2317_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0304_ : _0354_;
  assign _3208_ = _2318_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0004_ : _0066_;
  assign _3209_ = _2319_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0104_ : _0166_;
  assign _3210_ = _2320_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0204_ : _0266_;
  assign _3211_ = _2321_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0304_ : _0366_;
  assign _3212_ = _2322_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0004_ : _0078_;
  assign _3213_ = _2323_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0104_ : _0178_;
  assign _3214_ = _2324_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0204_ : _0278_;
  assign _3215_ = _2325_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0304_ : _0378_;
  assign _3216_ = _2326_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0004_ : _0090_;
  assign _3217_ = _2327_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0104_ : _0190_;
  assign _3218_ = _2328_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0204_ : _0290_;
  assign _3219_ = _2329_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3485" *) _0304_ : _0390_;
  assign _3220_ = _1527_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0004_ : _0005_;
  assign _3221_ = _1495_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3188_ : _3220_;
  assign _0406_ = _1463_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3156_ : _3221_;
  assign _3222_ = _1528_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0104_ : _0105_;
  assign _3223_ = _1496_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3189_ : _3222_;
  assign _0470_ = _1464_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3157_ : _3223_;
  assign _3224_ = _1529_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0204_ : _0205_;
  assign _3225_ = _1497_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3190_ : _3224_;
  assign _0534_ = _1465_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3158_ : _3225_;
  assign _3226_ = _1530_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0304_ : _0305_;
  assign _3227_ = _1498_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3191_ : _3226_;
  assign _0598_ = _1466_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3159_ : _3227_;
  assign _3228_ = _1531_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0004_ : _0018_;
  assign _3229_ = _1499_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3192_ : _3228_;
  assign _0414_ = _1467_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3160_ : _3229_;
  assign _3230_ = _1532_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0104_ : _0118_;
  assign _3231_ = _1500_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3193_ : _3230_;
  assign _0478_ = _1468_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3161_ : _3231_;
  assign _3232_ = _1533_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0204_ : _0218_;
  assign _3233_ = _1501_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3194_ : _3232_;
  assign _0542_ = _1469_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3162_ : _3233_;
  assign _3234_ = _1534_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0304_ : _0318_;
  assign _3235_ = _1502_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3195_ : _3234_;
  assign _0606_ = _1470_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3163_ : _3235_;
  assign _3236_ = _1535_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0004_ : _0030_;
  assign _3237_ = _1503_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3196_ : _3236_;
  assign _0422_ = _1471_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3164_ : _3237_;
  assign _3238_ = _1536_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0104_ : _0130_;
  assign _3239_ = _1504_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3197_ : _3238_;
  assign _0486_ = _1472_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3165_ : _3239_;
  assign _3240_ = _1537_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0204_ : _0230_;
  assign _3241_ = _1505_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3198_ : _3240_;
  assign _0550_ = _1473_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3166_ : _3241_;
  assign _3242_ = _1538_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0304_ : _0330_;
  assign _3243_ = _1506_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3199_ : _3242_;
  assign _0614_ = _1474_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3167_ : _3243_;
  assign _3244_ = _1539_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0004_ : _0042_;
  assign _3245_ = _1507_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3200_ : _3244_;
  assign _0430_ = _1475_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3168_ : _3245_;
  assign _3246_ = _1540_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0104_ : _0142_;
  assign _3247_ = _1508_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3201_ : _3246_;
  assign _0494_ = _1476_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3169_ : _3247_;
  assign _3248_ = _1541_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0204_ : _0242_;
  assign _3249_ = _1509_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3202_ : _3248_;
  assign _0558_ = _1477_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3170_ : _3249_;
  assign _3250_ = _1542_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0304_ : _0342_;
  assign _3251_ = _1510_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3203_ : _3250_;
  assign _0622_ = _1478_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3171_ : _3251_;
  assign _3252_ = _1543_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0004_ : _0054_;
  assign _3253_ = _1511_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3204_ : _3252_;
  assign _0438_ = _1479_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3172_ : _3253_;
  assign _3254_ = _1544_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0104_ : _0154_;
  assign _3255_ = _1512_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3205_ : _3254_;
  assign _0502_ = _1480_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3173_ : _3255_;
  assign _3256_ = _1545_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0204_ : _0254_;
  assign _3257_ = _1513_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3206_ : _3256_;
  assign _0566_ = _1481_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3174_ : _3257_;
  assign _3258_ = _1546_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0304_ : _0354_;
  assign _3259_ = _1514_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3207_ : _3258_;
  assign _0630_ = _1482_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3175_ : _3259_;
  assign _3260_ = _1547_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0004_ : _0066_;
  assign _3261_ = _1515_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3208_ : _3260_;
  assign _0446_ = _1483_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3176_ : _3261_;
  assign _3262_ = _1548_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0104_ : _0166_;
  assign _3263_ = _1516_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3209_ : _3262_;
  assign _0510_ = _1484_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3177_ : _3263_;
  assign _3264_ = _1549_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0204_ : _0266_;
  assign _3265_ = _1517_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3210_ : _3264_;
  assign _0574_ = _1485_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3178_ : _3265_;
  assign _3266_ = _1550_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0304_ : _0366_;
  assign _3267_ = _1518_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3211_ : _3266_;
  assign _0638_ = _1486_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3179_ : _3267_;
  assign _3268_ = _1551_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0004_ : _0078_;
  assign _3269_ = _1519_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3212_ : _3268_;
  assign _0454_ = _1487_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3180_ : _3269_;
  assign _3270_ = _1552_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0104_ : _0178_;
  assign _3271_ = _1520_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3213_ : _3270_;
  assign _0518_ = _1488_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3181_ : _3271_;
  assign _3272_ = _1553_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0204_ : _0278_;
  assign _3273_ = _1521_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3214_ : _3272_;
  assign _0582_ = _1489_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3182_ : _3273_;
  assign _3274_ = _1554_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0304_ : _0378_;
  assign _3275_ = _1522_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3215_ : _3274_;
  assign _0646_ = _1490_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3183_ : _3275_;
  assign _3276_ = _1555_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0004_ : _0090_;
  assign _3277_ = _1523_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3216_ : _3276_;
  assign _0462_ = _1491_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3184_ : _3277_;
  assign _3278_ = _1556_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0104_ : _0190_;
  assign _3279_ = _1524_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3217_ : _3278_;
  assign _0526_ = _1492_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3185_ : _3279_;
  assign _3280_ = _1557_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0204_ : _0290_;
  assign _3281_ = _1525_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3218_ : _3280_;
  assign _0590_ = _1493_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3186_ : _3281_;
  assign _3282_ = _1558_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _0304_ : _0390_;
  assign _3283_ = _1526_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3219_ : _3282_;
  assign _0654_ = _1494_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3486" *) _3187_ : _3283_;
  assign _3284_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0400_ : { _0404_, _0402_ };
  assign _0407_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0406_ : _3284_;
  assign _3285_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0464_ : { _0468_, _0466_ };
  assign _0471_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0470_ : _3285_;
  assign _3286_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0528_ : { _0532_, _0530_ };
  assign _0535_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0534_ : _3286_;
  assign _3287_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0592_ : { _0596_, _0594_ };
  assign _0599_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0598_ : _3287_;
  assign _3288_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0408_ : { _0412_, _0410_ };
  assign _0415_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0414_ : _3288_;
  assign _3289_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0472_ : { _0476_, _0474_ };
  assign _0479_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0478_ : _3289_;
  assign _3290_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0536_ : { _0540_, _0538_ };
  assign _0543_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0542_ : _3290_;
  assign _3291_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0600_ : { _0604_, _0602_ };
  assign _0607_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0606_ : _3291_;
  assign _3292_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0416_ : { _0420_, _0418_ };
  assign _0423_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0422_ : _3292_;
  assign _3293_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0480_ : { _0484_, _0482_ };
  assign _0487_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0486_ : _3293_;
  assign _3294_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0544_ : { _0548_, _0546_ };
  assign _0551_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0550_ : _3294_;
  assign _3295_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0608_ : { _0612_, _0610_ };
  assign _0615_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0614_ : _3295_;
  assign _3296_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0424_ : { _0428_, _0426_ };
  assign _0431_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0430_ : _3296_;
  assign _3297_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0488_ : { _0492_, _0490_ };
  assign _0495_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0494_ : _3297_;
  assign _3298_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0552_ : { _0556_, _0554_ };
  assign _0559_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0558_ : _3298_;
  assign _3299_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0616_ : { _0620_, _0618_ };
  assign _0623_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0622_ : _3299_;
  assign _3300_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0432_ : { _0436_, _0434_ };
  assign _0439_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0438_ : _3300_;
  assign _3301_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0496_ : { _0500_, _0498_ };
  assign _0503_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0502_ : _3301_;
  assign _3302_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0560_ : { _0564_, _0562_ };
  assign _0567_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0566_ : _3302_;
  assign _3303_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0624_ : { _0628_, _0626_ };
  assign _0631_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0630_ : _3303_;
  assign _3304_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0440_ : { _0444_, _0442_ };
  assign _0447_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0446_ : _3304_;
  assign _3305_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0504_ : { _0508_, _0506_ };
  assign _0511_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0510_ : _3305_;
  assign _3306_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0568_ : { _0572_, _0570_ };
  assign _0575_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0574_ : _3306_;
  assign _3307_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0632_ : { _0636_, _0634_ };
  assign _0639_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0638_ : _3307_;
  assign _3308_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0448_ : { _0452_, _0450_ };
  assign _0455_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0454_ : _3308_;
  assign _3309_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0512_ : { _0516_, _0514_ };
  assign _0519_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0518_ : _3309_;
  assign _3310_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0576_ : { _0580_, _0578_ };
  assign _0583_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0582_ : _3310_;
  assign _3311_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0640_ : { _0644_, _0642_ };
  assign _0647_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0646_ : _3311_;
  assign _3312_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0456_ : { _0460_, _0458_ };
  assign _0463_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0462_ : _3312_;
  assign _3313_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0520_ : { _0524_, _0522_ };
  assign _0527_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0526_ : _3313_;
  assign _3314_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0584_ : { _0588_, _0586_ };
  assign _0591_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0590_ : _3314_;
  assign _3315_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0648_ : { _0652_, _0650_ };
  assign _0655_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3488" *) _0654_ : _3315_;
  assign _0010_ = _1559_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0000_ : _0002_;
  assign _0110_ = _1560_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0100_ : _0102_;
  assign _0210_ = _1561_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0200_ : _0202_;
  assign _0310_ = _1562_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0300_ : _0302_;
  assign _0022_ = _1563_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0000_ : _0016_;
  assign _0122_ = _1564_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0100_ : _0116_;
  assign _0222_ = _1565_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0200_ : _0216_;
  assign _0322_ = _1566_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0300_ : _0316_;
  assign _0034_ = _1567_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0000_ : _0028_;
  assign _0134_ = _1568_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0100_ : _0128_;
  assign _0234_ = _1569_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0200_ : _0228_;
  assign _0334_ = _1570_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0300_ : _0328_;
  assign _0046_ = _1571_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0000_ : _0040_;
  assign _0146_ = _1572_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0100_ : _0140_;
  assign _0246_ = _1573_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0200_ : _0240_;
  assign _0346_ = _1574_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0300_ : _0340_;
  assign _0058_ = _1575_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0000_ : _0052_;
  assign _0158_ = _1576_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0100_ : _0152_;
  assign _0258_ = _1577_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0200_ : _0252_;
  assign _0358_ = _1578_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0300_ : _0352_;
  assign _0070_ = _1579_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0000_ : _0064_;
  assign _0170_ = _1580_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0100_ : _0164_;
  assign _0270_ = _1581_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0200_ : _0264_;
  assign _0370_ = _1582_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0300_ : _0364_;
  assign _0082_ = _1583_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0000_ : _0076_;
  assign _0182_ = _1584_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0100_ : _0176_;
  assign _0282_ = _1585_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0200_ : _0276_;
  assign _0382_ = _1586_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0300_ : _0376_;
  assign _0094_ = _1587_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0000_ : _0088_;
  assign _0194_ = _1588_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0100_ : _0188_;
  assign _0294_ = _1589_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0200_ : _0288_;
  assign _0394_ = _1590_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3523" *) _0300_ : _0388_;
  assign _0012_ = _1591_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0001_ : _0003_;
  assign _0112_ = _1592_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0101_ : _0103_;
  assign _0212_ = _1593_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0201_ : _0203_;
  assign _0312_ = _1594_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0301_ : _0303_;
  assign _0024_ = _1595_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0001_ : _0017_;
  assign _0124_ = _1596_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0101_ : _0117_;
  assign _0224_ = _1597_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0201_ : _0217_;
  assign _0324_ = _1598_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0301_ : _0317_;
  assign _0036_ = _1599_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0001_ : _0029_;
  assign _0136_ = _1600_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0101_ : _0129_;
  assign _0236_ = _1601_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0201_ : _0229_;
  assign _0336_ = _1602_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0301_ : _0329_;
  assign _0048_ = _1603_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0001_ : _0041_;
  assign _0148_ = _1604_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0101_ : _0141_;
  assign _0248_ = _1605_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0201_ : _0241_;
  assign _0348_ = _1606_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0301_ : _0341_;
  assign _0060_ = _1607_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0001_ : _0053_;
  assign _0160_ = _1608_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0101_ : _0153_;
  assign _0260_ = _1609_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0201_ : _0253_;
  assign _0360_ = _1610_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0301_ : _0353_;
  assign _0072_ = _1611_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0001_ : _0065_;
  assign _0172_ = _1612_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0101_ : _0165_;
  assign _0272_ = _1613_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0201_ : _0265_;
  assign _0372_ = _1614_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0301_ : _0365_;
  assign _0084_ = _1615_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0001_ : _0077_;
  assign _0184_ = _1616_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0101_ : _0177_;
  assign _0284_ = _1617_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0201_ : _0277_;
  assign _0384_ = _1618_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0301_ : _0377_;
  assign _0096_ = _1619_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0001_ : _0089_;
  assign _0196_ = _1620_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0101_ : _0189_;
  assign _0296_ = _1621_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0201_ : _0289_;
  assign _0396_ = _1622_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3524" *) _0301_ : _0389_;
  assign _0008_ = _1623_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0006_ : _0007_;
  assign _0108_ = _1624_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0106_ : _0107_;
  assign _0208_ = _1625_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0206_ : _0207_;
  assign _0308_ = _1626_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0306_ : _0307_;
  assign _0020_ = _1627_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0006_ : _0019_;
  assign _0120_ = _1628_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0106_ : _0119_;
  assign _0220_ = _1629_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0206_ : _0219_;
  assign _0320_ = _1630_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0306_ : _0319_;
  assign _0032_ = _1631_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0006_ : _0031_;
  assign _0132_ = _1632_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0106_ : _0131_;
  assign _0232_ = _1633_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0206_ : _0231_;
  assign _0332_ = _1634_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0306_ : _0331_;
  assign _0044_ = _1635_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0006_ : _0043_;
  assign _0144_ = _1636_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0106_ : _0143_;
  assign _0244_ = _1637_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0206_ : _0243_;
  assign _0344_ = _1638_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0306_ : _0343_;
  assign _0056_ = _1639_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0006_ : _0055_;
  assign _0156_ = _1640_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0106_ : _0155_;
  assign _0256_ = _1641_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0206_ : _0255_;
  assign _0356_ = _1642_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0306_ : _0355_;
  assign _0068_ = _1643_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0006_ : _0067_;
  assign _0168_ = _1644_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0106_ : _0167_;
  assign _0268_ = _1645_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0206_ : _0267_;
  assign _0368_ = _1646_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0306_ : _0367_;
  assign _0080_ = _1647_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0006_ : _0079_;
  assign _0180_ = _1648_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0106_ : _0179_;
  assign _0280_ = _1649_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0206_ : _0279_;
  assign _0380_ = _1650_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0306_ : _0379_;
  assign _0092_ = _1651_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0006_ : _0091_;
  assign _0192_ = _1652_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0106_ : _0191_;
  assign _0292_ = _1653_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0206_ : _0291_;
  assign _0392_ = _1654_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3525" *) _0306_ : _0391_;
  assign _3316_ = _1527_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0005_ : _0004_;
  assign _3317_ = _1495_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3156_ : _3316_;
  assign _0014_ = _1463_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3188_ : _3317_;
  assign _3318_ = _1528_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0105_ : _0104_;
  assign _3319_ = _1496_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3157_ : _3318_;
  assign _0114_ = _1464_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3189_ : _3319_;
  assign _3320_ = _1529_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0205_ : _0204_;
  assign _3321_ = _1497_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3158_ : _3320_;
  assign _0214_ = _1465_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3190_ : _3321_;
  assign _3322_ = _1530_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0305_ : _0304_;
  assign _3323_ = _1498_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3159_ : _3322_;
  assign _0314_ = _1466_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3191_ : _3323_;
  assign _3324_ = _1531_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0018_ : _0004_;
  assign _3325_ = _1499_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3160_ : _3324_;
  assign _0026_ = _1467_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3192_ : _3325_;
  assign _3326_ = _1532_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0118_ : _0104_;
  assign _3327_ = _1500_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3161_ : _3326_;
  assign _0126_ = _1468_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3193_ : _3327_;
  assign _3328_ = _1533_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0218_ : _0204_;
  assign _3329_ = _1501_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3162_ : _3328_;
  assign _0226_ = _1469_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3194_ : _3329_;
  assign _3330_ = _1534_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0318_ : _0304_;
  assign _3331_ = _1502_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3163_ : _3330_;
  assign _0326_ = _1470_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3195_ : _3331_;
  assign _3332_ = _1535_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0030_ : _0004_;
  assign _3333_ = _1503_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3164_ : _3332_;
  assign _0038_ = _1471_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3196_ : _3333_;
  assign _3334_ = _1536_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0130_ : _0104_;
  assign _3335_ = _1504_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3165_ : _3334_;
  assign _0138_ = _1472_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3197_ : _3335_;
  assign _3336_ = _1537_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0230_ : _0204_;
  assign _3337_ = _1505_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3166_ : _3336_;
  assign _0238_ = _1473_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3198_ : _3337_;
  assign _3338_ = _1538_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0330_ : _0304_;
  assign _3339_ = _1506_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3167_ : _3338_;
  assign _0338_ = _1474_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3199_ : _3339_;
  assign _3340_ = _1539_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0042_ : _0004_;
  assign _3341_ = _1507_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3168_ : _3340_;
  assign _0050_ = _1475_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3200_ : _3341_;
  assign _3342_ = _1540_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0142_ : _0104_;
  assign _3343_ = _1508_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3169_ : _3342_;
  assign _0150_ = _1476_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3201_ : _3343_;
  assign _3344_ = _1541_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0242_ : _0204_;
  assign _3345_ = _1509_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3170_ : _3344_;
  assign _0250_ = _1477_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3202_ : _3345_;
  assign _3346_ = _1542_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0342_ : _0304_;
  assign _3347_ = _1510_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3171_ : _3346_;
  assign _0350_ = _1478_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3203_ : _3347_;
  assign _3348_ = _1543_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0054_ : _0004_;
  assign _3349_ = _1511_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3172_ : _3348_;
  assign _0062_ = _1479_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3204_ : _3349_;
  assign _3350_ = _1544_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0154_ : _0104_;
  assign _3351_ = _1512_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3173_ : _3350_;
  assign _0162_ = _1480_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3205_ : _3351_;
  assign _3352_ = _1545_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0254_ : _0204_;
  assign _3353_ = _1513_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3174_ : _3352_;
  assign _0262_ = _1481_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3206_ : _3353_;
  assign _3354_ = _1546_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0354_ : _0304_;
  assign _3355_ = _1514_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3175_ : _3354_;
  assign _0362_ = _1482_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3207_ : _3355_;
  assign _3356_ = _1547_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0066_ : _0004_;
  assign _3357_ = _1515_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3176_ : _3356_;
  assign _0074_ = _1483_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3208_ : _3357_;
  assign _3358_ = _1548_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0166_ : _0104_;
  assign _3359_ = _1516_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3177_ : _3358_;
  assign _0174_ = _1484_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3209_ : _3359_;
  assign _3360_ = _1549_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0266_ : _0204_;
  assign _3361_ = _1517_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3178_ : _3360_;
  assign _0274_ = _1485_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3210_ : _3361_;
  assign _3362_ = _1550_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0366_ : _0304_;
  assign _3363_ = _1518_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3179_ : _3362_;
  assign _0374_ = _1486_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3211_ : _3363_;
  assign _3364_ = _1551_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0078_ : _0004_;
  assign _3365_ = _1519_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3180_ : _3364_;
  assign _0086_ = _1487_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3212_ : _3365_;
  assign _3366_ = _1552_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0178_ : _0104_;
  assign _3367_ = _1520_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3181_ : _3366_;
  assign _0186_ = _1488_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3213_ : _3367_;
  assign _3368_ = _1553_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0278_ : _0204_;
  assign _3369_ = _1521_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3182_ : _3368_;
  assign _0286_ = _1489_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3214_ : _3369_;
  assign _3370_ = _1554_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0378_ : _0304_;
  assign _3371_ = _1522_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3183_ : _3370_;
  assign _0386_ = _1490_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3215_ : _3371_;
  assign _3372_ = _1555_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0090_ : _0004_;
  assign _3373_ = _1523_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3184_ : _3372_;
  assign _0098_ = _1491_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3216_ : _3373_;
  assign _3374_ = _1556_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0190_ : _0104_;
  assign _3375_ = _1524_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3185_ : _3374_;
  assign _0198_ = _1492_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3217_ : _3375_;
  assign _3376_ = _1557_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0290_ : _0204_;
  assign _3377_ = _1525_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3186_ : _3376_;
  assign _0298_ = _1493_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3218_ : _3377_;
  assign _3378_ = _1558_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _0390_ : _0304_;
  assign _3379_ = _1526_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3187_ : _3378_;
  assign _0398_ = _1494_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3528" *) _3219_ : _3379_;
  assign _3380_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0008_ : { _0012_, _0010_ };
  assign _0015_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0014_ : _3380_;
  assign _3381_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0108_ : { _0112_, _0110_ };
  assign _0115_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0114_ : _3381_;
  assign _3382_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0208_ : { _0212_, _0210_ };
  assign _0215_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0214_ : _3382_;
  assign _3383_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0308_ : { _0312_, _0310_ };
  assign _0315_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0314_ : _3383_;
  assign _3384_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0020_ : { _0024_, _0022_ };
  assign _0027_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0026_ : _3384_;
  assign _3385_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0120_ : { _0124_, _0122_ };
  assign _0127_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0126_ : _3385_;
  assign _3386_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0220_ : { _0224_, _0222_ };
  assign _0227_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0226_ : _3386_;
  assign _3387_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0320_ : { _0324_, _0322_ };
  assign _0327_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0326_ : _3387_;
  assign _3388_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0032_ : { _0036_, _0034_ };
  assign _0039_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0038_ : _3388_;
  assign _3389_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0132_ : { _0136_, _0134_ };
  assign _0139_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0138_ : _3389_;
  assign _3390_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0232_ : { _0236_, _0234_ };
  assign _0239_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0238_ : _3390_;
  assign _3391_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0332_ : { _0336_, _0334_ };
  assign _0339_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0338_ : _3391_;
  assign _3392_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0044_ : { _0048_, _0046_ };
  assign _0051_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0050_ : _3392_;
  assign _3393_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0144_ : { _0148_, _0146_ };
  assign _0151_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0150_ : _3393_;
  assign _3394_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0244_ : { _0248_, _0246_ };
  assign _0251_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0250_ : _3394_;
  assign _3395_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0344_ : { _0348_, _0346_ };
  assign _0351_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0350_ : _3395_;
  assign _3396_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0056_ : { _0060_, _0058_ };
  assign _0063_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0062_ : _3396_;
  assign _3397_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0156_ : { _0160_, _0158_ };
  assign _0163_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0162_ : _3397_;
  assign _3398_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0256_ : { _0260_, _0258_ };
  assign _0263_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0262_ : _3398_;
  assign _3399_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0356_ : { _0360_, _0358_ };
  assign _0363_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0362_ : _3399_;
  assign _3400_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0068_ : { _0072_, _0070_ };
  assign _0075_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0074_ : _3400_;
  assign _3401_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0168_ : { _0172_, _0170_ };
  assign _0175_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0174_ : _3401_;
  assign _3402_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0268_ : { _0272_, _0270_ };
  assign _0275_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0274_ : _3402_;
  assign _3403_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0368_ : { _0372_, _0370_ };
  assign _0375_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0374_ : _3403_;
  assign _3404_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0080_ : { _0084_, _0082_ };
  assign _0087_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0086_ : _3404_;
  assign _3405_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0180_ : { _0184_, _0182_ };
  assign _0187_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0186_ : _3405_;
  assign _3406_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0280_ : { _0284_, _0282_ };
  assign _0287_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0286_ : _3406_;
  assign _3407_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0380_ : { _0384_, _0382_ };
  assign _0387_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0386_ : _3407_;
  assign _3408_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0092_ : { _0096_, _0094_ };
  assign _0099_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0098_ : _3408_;
  assign _3409_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0192_ : { _0196_, _0194_ };
  assign _0199_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0198_ : _3409_;
  assign _3410_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0292_ : { _0296_, _0294_ };
  assign _0299_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0298_ : _3410_;
  assign _3411_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0392_ : { _0396_, _0394_ };
  assign _0399_ = reg2dp_fp16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3530" *) _0398_ : _3411_;
  assign { _0657_, _0656_ } = _1655_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign { _0737_, _0736_ } = _1655_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign { _0817_, _0816_ } = _1655_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign { _0897_, _0896_ } = _1655_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign { _0667_, _0666_ } = _1656_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign { _0747_, _0746_ } = _1656_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign { _0827_, _0826_ } = _1656_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign { _0907_, _0906_ } = _1656_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign { _0677_, _0676_ } = _1657_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign { _0757_, _0756_ } = _1657_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign { _0837_, _0836_ } = _1657_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign { _0917_, _0916_ } = _1657_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign { _0687_, _0686_ } = _1658_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign { _0767_, _0766_ } = _1658_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign { _0847_, _0846_ } = _1658_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign { _0927_, _0926_ } = _1658_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign { _0697_, _0696_ } = _1659_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign { _0777_, _0776_ } = _1659_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign { _0857_, _0856_ } = _1659_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign { _0937_, _0936_ } = _1659_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign { _0707_, _0706_ } = _1660_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign { _0787_, _0786_ } = _1660_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign { _0867_, _0866_ } = _1660_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign { _0947_, _0946_ } = _1660_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign { _0717_, _0716_ } = _1661_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign { _0797_, _0796_ } = _1661_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign { _0877_, _0876_ } = _1661_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign { _0957_, _0956_ } = _1661_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign { _0727_, _0726_ } = _1662_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign { _0807_, _0806_ } = _1662_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign { _0887_, _0886_ } = _1662_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign { _0967_, _0966_ } = _1662_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3552" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign { _0659_, _0658_ } = _1655_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data0[27:0] : 28'b0000000000000000000000000000;
  assign { _0739_, _0738_ } = _1655_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data0[55:28] : 28'b0000000000000000000000000000;
  assign { _0819_, _0818_ } = _1655_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data0[83:56] : 28'b0000000000000000000000000000;
  assign { _0899_, _0898_ } = _1655_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data0[111:84] : 28'b0000000000000000000000000000;
  assign { _0669_, _0668_ } = _1656_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data1[27:0] : 28'b0000000000000000000000000000;
  assign { _0749_, _0748_ } = _1656_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data1[55:28] : 28'b0000000000000000000000000000;
  assign { _0829_, _0828_ } = _1656_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data1[83:56] : 28'b0000000000000000000000000000;
  assign { _0909_, _0908_ } = _1656_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data1[111:84] : 28'b0000000000000000000000000000;
  assign { _0679_, _0678_ } = _1657_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data2[27:0] : 28'b0000000000000000000000000000;
  assign { _0759_, _0758_ } = _1657_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data2[55:28] : 28'b0000000000000000000000000000;
  assign { _0839_, _0838_ } = _1657_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data2[83:56] : 28'b0000000000000000000000000000;
  assign { _0919_, _0918_ } = _1657_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data2[111:84] : 28'b0000000000000000000000000000;
  assign { _0689_, _0688_ } = _1658_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data3[27:0] : 28'b0000000000000000000000000000;
  assign { _0769_, _0768_ } = _1658_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data3[55:28] : 28'b0000000000000000000000000000;
  assign { _0849_, _0848_ } = _1658_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data3[83:56] : 28'b0000000000000000000000000000;
  assign { _0929_, _0928_ } = _1658_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data3[111:84] : 28'b0000000000000000000000000000;
  assign { _0699_, _0698_ } = _1659_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data4[27:0] : 28'b0000000000000000000000000000;
  assign { _0779_, _0778_ } = _1659_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data4[55:28] : 28'b0000000000000000000000000000;
  assign { _0859_, _0858_ } = _1659_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data4[83:56] : 28'b0000000000000000000000000000;
  assign { _0939_, _0938_ } = _1659_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data4[111:84] : 28'b0000000000000000000000000000;
  assign { _0709_, _0708_ } = _1660_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data5[27:0] : 28'b0000000000000000000000000000;
  assign { _0789_, _0788_ } = _1660_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data5[55:28] : 28'b0000000000000000000000000000;
  assign { _0869_, _0868_ } = _1660_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data5[83:56] : 28'b0000000000000000000000000000;
  assign { _0949_, _0948_ } = _1660_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data5[111:84] : 28'b0000000000000000000000000000;
  assign { _0719_, _0718_ } = _1661_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data6[27:0] : 28'b0000000000000000000000000000;
  assign { _0799_, _0798_ } = _1661_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data6[55:28] : 28'b0000000000000000000000000000;
  assign { _0879_, _0878_ } = _1661_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data6[83:56] : 28'b0000000000000000000000000000;
  assign { _0959_, _0958_ } = _1661_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data6[111:84] : 28'b0000000000000000000000000000;
  assign { _0729_, _0728_ } = _1662_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data7[27:0] : 28'b0000000000000000000000000000;
  assign { _0809_, _0808_ } = _1662_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data7[55:28] : 28'b0000000000000000000000000000;
  assign { _0889_, _0888_ } = _1662_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data7[83:56] : 28'b0000000000000000000000000000;
  assign { _0969_, _0968_ } = _1662_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3553" *) mem_data7[111:84] : 28'b0000000000000000000000000000;
  assign _0660_ = _1663_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign _0740_ = _1663_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign _0820_ = _1663_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign _0900_ = _1663_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign _0670_ = _1664_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign _0750_ = _1664_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign _0830_ = _1664_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign _0910_ = _1664_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign _0680_ = _1665_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign _0760_ = _1665_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign _0840_ = _1665_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign _0920_ = _1665_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign _0690_ = _1666_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign _0770_ = _1666_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign _0850_ = _1666_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign _0930_ = _1666_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign _0700_ = _1667_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign _0780_ = _1667_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign _0860_ = _1667_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign _0940_ = _1667_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign _0710_ = _1668_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign _0790_ = _1668_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign _0870_ = _1668_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign _0950_ = _1668_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign _0720_ = _1669_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign _0800_ = _1669_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign _0880_ = _1669_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign _0960_ = _1669_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign _0730_ = _1670_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[27:0] : 28'b0000000000000000000000000000;
  assign _0810_ = _1670_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[55:28] : 28'b0000000000000000000000000000;
  assign _0890_ = _1670_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[83:56] : 28'b0000000000000000000000000000;
  assign _0970_ = _1670_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3554" *) datin_buf_2d[111:84] : 28'b0000000000000000000000000000;
  assign _0661_ = _1663_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data0[27:0] : 28'b0000000000000000000000000000;
  assign _0741_ = _1663_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data0[55:28] : 28'b0000000000000000000000000000;
  assign _0821_ = _1663_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data0[83:56] : 28'b0000000000000000000000000000;
  assign _0901_ = _1663_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data0[111:84] : 28'b0000000000000000000000000000;
  assign _0671_ = _1664_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data1[27:0] : 28'b0000000000000000000000000000;
  assign _0751_ = _1664_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data1[55:28] : 28'b0000000000000000000000000000;
  assign _0831_ = _1664_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data1[83:56] : 28'b0000000000000000000000000000;
  assign _0911_ = _1664_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data1[111:84] : 28'b0000000000000000000000000000;
  assign _0681_ = _1665_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data2[27:0] : 28'b0000000000000000000000000000;
  assign _0761_ = _1665_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data2[55:28] : 28'b0000000000000000000000000000;
  assign _0841_ = _1665_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data2[83:56] : 28'b0000000000000000000000000000;
  assign _0921_ = _1665_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data2[111:84] : 28'b0000000000000000000000000000;
  assign _0691_ = _1666_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data3[27:0] : 28'b0000000000000000000000000000;
  assign _0771_ = _1666_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data3[55:28] : 28'b0000000000000000000000000000;
  assign _0851_ = _1666_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data3[83:56] : 28'b0000000000000000000000000000;
  assign _0931_ = _1666_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data3[111:84] : 28'b0000000000000000000000000000;
  assign _0701_ = _1667_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data4[27:0] : 28'b0000000000000000000000000000;
  assign _0781_ = _1667_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data4[55:28] : 28'b0000000000000000000000000000;
  assign _0861_ = _1667_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data4[83:56] : 28'b0000000000000000000000000000;
  assign _0941_ = _1667_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data4[111:84] : 28'b0000000000000000000000000000;
  assign _0711_ = _1668_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data5[27:0] : 28'b0000000000000000000000000000;
  assign _0791_ = _1668_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data5[55:28] : 28'b0000000000000000000000000000;
  assign _0871_ = _1668_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data5[83:56] : 28'b0000000000000000000000000000;
  assign _0951_ = _1668_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data5[111:84] : 28'b0000000000000000000000000000;
  assign _0721_ = _1669_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data6[27:0] : 28'b0000000000000000000000000000;
  assign _0801_ = _1669_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data6[55:28] : 28'b0000000000000000000000000000;
  assign _0881_ = _1669_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data6[83:56] : 28'b0000000000000000000000000000;
  assign _0961_ = _1669_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data6[111:84] : 28'b0000000000000000000000000000;
  assign _0731_ = _1670_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data7[27:0] : 28'b0000000000000000000000000000;
  assign _0811_ = _1670_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data7[55:28] : 28'b0000000000000000000000000000;
  assign _0891_ = _1670_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data7[83:56] : 28'b0000000000000000000000000000;
  assign _0971_ = _1670_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3555" *) mem_data7[111:84] : 28'b0000000000000000000000000000;
  assign _0662_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0663_ : { _0665_, _0664_ };
  assign _0742_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0743_ : { _0745_, _0744_ };
  assign _0822_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0823_ : { _0825_, _0824_ };
  assign _0902_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0903_ : { _0905_, _0904_ };
  assign _0672_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0673_ : { _0675_, _0674_ };
  assign _0752_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0753_ : { _0755_, _0754_ };
  assign _0832_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0833_ : { _0835_, _0834_ };
  assign _0912_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0913_ : { _0915_, _0914_ };
  assign _0682_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0683_ : { _0685_, _0684_ };
  assign _0762_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0763_ : { _0765_, _0764_ };
  assign _0842_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0843_ : { _0845_, _0844_ };
  assign _0922_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0923_ : { _0925_, _0924_ };
  assign _0692_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0693_ : { _0695_, _0694_ };
  assign _0772_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0773_ : { _0775_, _0774_ };
  assign _0852_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0853_ : { _0855_, _0854_ };
  assign _0932_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0933_ : { _0935_, _0934_ };
  assign _0702_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0703_ : { _0705_, _0704_ };
  assign _0782_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0783_ : { _0785_, _0784_ };
  assign _0862_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0863_ : { _0865_, _0864_ };
  assign _0942_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0943_ : { _0945_, _0944_ };
  assign _0712_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0713_ : { _0715_, _0714_ };
  assign _0792_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0793_ : { _0795_, _0794_ };
  assign _0872_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0873_ : { _0875_, _0874_ };
  assign _0952_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0953_ : { _0955_, _0954_ };
  assign _0722_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0723_ : { _0725_, _0724_ };
  assign _0802_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0803_ : { _0805_, _0804_ };
  assign _0882_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0883_ : { _0885_, _0884_ };
  assign _0962_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0963_ : { _0965_, _0964_ };
  assign _0732_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0733_ : { _0735_, _0734_ };
  assign _0812_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0813_ : { _0815_, _0814_ };
  assign _0892_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0893_ : { _0895_, _0894_ };
  assign _0972_ = reg2dp_int16_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3564" *) _0973_ : { _0975_, _0974_ };
  assign _3412_ = _0977_[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) datin_buf_2d[27:0] : mem_data0[27:0];
  assign _1932_[27:0] = _2638_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0407_ : _3412_;
  assign _3413_ = _0977_[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) datin_buf_2d[27:0] : mem_data1[27:0];
  assign _1933_[27:0] = _2639_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0415_ : _3413_;
  assign _3414_ = _0977_[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) datin_buf_2d[27:0] : mem_data2[27:0];
  assign _1934_[27:0] = _2640_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0423_ : _3414_;
  assign _3415_ = _0977_[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) datin_buf_2d[27:0] : mem_data3[27:0];
  assign _1935_[27:0] = _2641_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0431_ : _3415_;
  assign _3416_ = _0977_[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) datin_buf_2d[27:0] : mem_data4[27:0];
  assign _1936_[27:0] = _2642_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0439_ : _3416_;
  assign _3417_ = _0977_[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) datin_buf_2d[27:0] : mem_data5[27:0];
  assign _1937_[27:0] = _2643_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0447_ : _3417_;
  assign _3418_ = _0977_[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) datin_buf_2d[27:0] : mem_data6[27:0];
  assign _1938_[27:0] = _2644_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0455_ : _3418_;
  assign _3419_ = _0977_[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) datin_buf_2d[27:0] : mem_data7[27:0];
  assign _1939_[27:0] = _2645_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3596" *) _0463_ : _3419_;
  assign _1940_[27:0] = _2638_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0015_ : _3412_;
  assign _3420_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1940_[27:0] : 28'b0000000000000000000000000000;
  assign _3421_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1932_[27:0] : _3420_[27:0];
  assign _0976_[27:0] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0662_ : _3421_[27:0];
  assign _1941_[27:0] = _2639_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0027_ : _3413_;
  assign _3422_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1941_[27:0] : 28'b0000000000000000000000000000;
  assign _3423_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1933_[27:0] : _3422_[27:0];
  assign _0982_[27:0] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0672_ : _3423_[27:0];
  assign _1942_[27:0] = _2640_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0039_ : _3414_;
  assign _3424_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1942_[27:0] : 28'b0000000000000000000000000000;
  assign _3425_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1934_[27:0] : _3424_[27:0];
  assign _0985_[27:0] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0682_ : _3425_[27:0];
  assign _1943_[27:0] = _2641_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0051_ : _3415_;
  assign _3426_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1943_[27:0] : 28'b0000000000000000000000000000;
  assign _3427_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1935_[27:0] : _3426_[27:0];
  assign _0988_[27:0] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0692_ : _3427_[27:0];
  assign _1944_[27:0] = _2642_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0063_ : _3416_;
  assign _3428_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1944_[27:0] : 28'b0000000000000000000000000000;
  assign _3429_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1936_[27:0] : _3428_[27:0];
  assign _0991_[27:0] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0702_ : _3429_[27:0];
  assign _1945_[27:0] = _2643_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0075_ : _3417_;
  assign _3430_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1945_[27:0] : 28'b0000000000000000000000000000;
  assign _3431_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1937_[27:0] : _3430_[27:0];
  assign _0994_[27:0] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0712_ : _3431_[27:0];
  assign _1946_[27:0] = _2644_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0087_ : _3418_;
  assign _3432_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1946_[27:0] : 28'b0000000000000000000000000000;
  assign _3433_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1938_[27:0] : _3432_[27:0];
  assign _0997_[27:0] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0722_ : _3433_[27:0];
  assign _1947_[27:0] = _2645_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0099_ : _3419_;
  assign _3434_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1947_[27:0] : 28'b0000000000000000000000000000;
  assign _3435_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _1939_[27:0] : _3434_[27:0];
  assign _1000_[27:0] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3597" *) _0732_ : _3435_[27:0];
  assign _3436_ = _0977_[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) datin_buf_2d[55:28] : mem_data0[55:28];
  assign _1948_[27:0] = _2646_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0471_ : _3436_;
  assign _3437_ = _0977_[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) datin_buf_2d[55:28] : mem_data1[55:28];
  assign _1949_[27:0] = _2647_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0479_ : _3437_;
  assign _3438_ = _0977_[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) datin_buf_2d[55:28] : mem_data2[55:28];
  assign _1950_[27:0] = _2648_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0487_ : _3438_;
  assign _3439_ = _0977_[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) datin_buf_2d[55:28] : mem_data3[55:28];
  assign _1951_[27:0] = _2649_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0495_ : _3439_;
  assign _3440_ = _0977_[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) datin_buf_2d[55:28] : mem_data4[55:28];
  assign _1952_[27:0] = _2650_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0503_ : _3440_;
  assign _3441_ = _0977_[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) datin_buf_2d[55:28] : mem_data5[55:28];
  assign _1953_[27:0] = _2651_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0511_ : _3441_;
  assign _3442_ = _0977_[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) datin_buf_2d[55:28] : mem_data6[55:28];
  assign _1954_[27:0] = _2652_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0519_ : _3442_;
  assign _3443_ = _0977_[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) datin_buf_2d[55:28] : mem_data7[55:28];
  assign _1955_[27:0] = _2653_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3599" *) _0527_ : _3443_;
  assign _1956_[27:0] = _2646_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0115_ : _3436_;
  assign _1957_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1956_[27:0] : 28'b0000000000000000000000000000;
  assign _3444_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1948_[27:0] : _1957_[27:0];
  assign _0976_[55:28] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0742_ : _3444_[27:0];
  assign _1958_[27:0] = _2647_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0127_ : _3437_;
  assign _3445_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1958_[27:0] : 28'b0000000000000000000000000000;
  assign _3446_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1949_[27:0] : _3445_[27:0];
  assign _0982_[55:28] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0752_ : _3446_[27:0];
  assign _1959_[27:0] = _2648_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0139_ : _3438_;
  assign _3447_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1959_[27:0] : 28'b0000000000000000000000000000;
  assign _3448_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1950_[27:0] : _3447_[27:0];
  assign _0985_[55:28] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0762_ : _3448_[27:0];
  assign _1960_[27:0] = _2649_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0151_ : _3439_;
  assign _3449_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1960_[27:0] : 28'b0000000000000000000000000000;
  assign _3450_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1951_[27:0] : _3449_[27:0];
  assign _0988_[55:28] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0772_ : _3450_[27:0];
  assign _1961_[27:0] = _2650_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0163_ : _3440_;
  assign _3451_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1961_[27:0] : 28'b0000000000000000000000000000;
  assign _3452_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1952_[27:0] : _3451_[27:0];
  assign _0991_[55:28] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0782_ : _3452_[27:0];
  assign _1962_[27:0] = _2651_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0175_ : _3441_;
  assign _3453_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1962_[27:0] : 28'b0000000000000000000000000000;
  assign _3454_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1953_[27:0] : _3453_[27:0];
  assign _0994_[55:28] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0792_ : _3454_[27:0];
  assign _1963_[27:0] = _2652_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0187_ : _3442_;
  assign _3455_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1963_[27:0] : 28'b0000000000000000000000000000;
  assign _3456_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1954_[27:0] : _3455_[27:0];
  assign _0997_[55:28] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0802_ : _3456_[27:0];
  assign _1964_[27:0] = _2653_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0199_ : _3443_;
  assign _3457_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1964_[27:0] : 28'b0000000000000000000000000000;
  assign _3458_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _1955_[27:0] : _3457_[27:0];
  assign _1000_[55:28] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3600" *) _0812_ : _3458_[27:0];
  assign _3459_ = _0977_[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) datin_buf_2d[83:56] : mem_data0[83:56];
  assign _1965_[27:0] = _2654_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0535_ : _3459_;
  assign _3460_ = _0977_[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) datin_buf_2d[83:56] : mem_data1[83:56];
  assign _1966_[27:0] = _2655_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0543_ : _3460_;
  assign _3461_ = _0977_[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) datin_buf_2d[83:56] : mem_data2[83:56];
  assign _1967_[27:0] = _2656_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0551_ : _3461_;
  assign _3462_ = _0977_[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) datin_buf_2d[83:56] : mem_data3[83:56];
  assign _1968_[27:0] = _2657_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0559_ : _3462_;
  assign _3463_ = _0977_[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) datin_buf_2d[83:56] : mem_data4[83:56];
  assign _1969_[27:0] = _2658_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0567_ : _3463_;
  assign _3464_ = _0977_[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) datin_buf_2d[83:56] : mem_data5[83:56];
  assign _1970_[27:0] = _2659_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0575_ : _3464_;
  assign _3465_ = _0977_[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) datin_buf_2d[83:56] : mem_data6[83:56];
  assign _1971_[27:0] = _2660_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0583_ : _3465_;
  assign _3466_ = _0977_[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) datin_buf_2d[83:56] : mem_data7[83:56];
  assign _1972_[27:0] = _2661_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3602" *) _0591_ : _3466_;
  assign _1973_[27:0] = _2654_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0215_ : _3459_;
  assign _3467_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1973_[27:0] : 28'b0000000000000000000000000000;
  assign _3468_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1965_[27:0] : _3467_[27:0];
  assign _0976_[83:56] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0822_ : _3468_[27:0];
  assign _1974_[27:0] = _2655_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0227_ : _3460_;
  assign _3469_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1974_[27:0] : 28'b0000000000000000000000000000;
  assign _3470_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1966_[27:0] : _3469_[27:0];
  assign _0982_[83:56] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0832_ : _3470_[27:0];
  assign _1975_[27:0] = _2656_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0239_ : _3461_;
  assign _3471_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1975_[27:0] : 28'b0000000000000000000000000000;
  assign _3472_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1967_[27:0] : _3471_[27:0];
  assign _0985_[83:56] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0842_ : _3472_[27:0];
  assign _1976_[27:0] = _2657_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0251_ : _3462_;
  assign _3473_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1976_[27:0] : 28'b0000000000000000000000000000;
  assign _3474_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1968_[27:0] : _3473_[27:0];
  assign _0988_[83:56] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0852_ : _3474_[27:0];
  assign _1977_[27:0] = _2658_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0263_ : _3463_;
  assign _3475_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1977_[27:0] : 28'b0000000000000000000000000000;
  assign _3476_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1969_[27:0] : _3475_[27:0];
  assign _0991_[83:56] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0862_ : _3476_[27:0];
  assign _1978_[27:0] = _2659_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0275_ : _3464_;
  assign _3477_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1978_[27:0] : 28'b0000000000000000000000000000;
  assign _3478_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1970_[27:0] : _3477_[27:0];
  assign _0994_[83:56] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0872_ : _3478_[27:0];
  assign _1979_[27:0] = _2660_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0287_ : _3465_;
  assign _3479_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1979_[27:0] : 28'b0000000000000000000000000000;
  assign _3480_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1971_[27:0] : _3479_[27:0];
  assign _0997_[83:56] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0882_ : _3480_[27:0];
  assign _1980_[27:0] = _2661_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0299_ : _3466_;
  assign _3481_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1980_[27:0] : 28'b0000000000000000000000000000;
  assign _3482_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _1972_[27:0] : _3481_[27:0];
  assign _1000_[83:56] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3603" *) _0892_ : _3482_[27:0];
  assign _3483_ = _0977_[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) datin_buf_2d[111:84] : mem_data0[111:84];
  assign _1981_[27:0] = _2662_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0599_ : _3483_;
  assign _3484_ = _0977_[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) datin_buf_2d[111:84] : mem_data1[111:84];
  assign _1982_[27:0] = _2663_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0607_ : _3484_;
  assign _3485_ = _0977_[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) datin_buf_2d[111:84] : mem_data2[111:84];
  assign _1983_[27:0] = _2664_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0615_ : _3485_;
  assign _3486_ = _0977_[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) datin_buf_2d[111:84] : mem_data3[111:84];
  assign _1984_[27:0] = _2665_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0623_ : _3486_;
  assign _3487_ = _0977_[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) datin_buf_2d[111:84] : mem_data4[111:84];
  assign _1985_[27:0] = _2666_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0631_ : _3487_;
  assign _3488_ = _0977_[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) datin_buf_2d[111:84] : mem_data5[111:84];
  assign _1986_[27:0] = _2667_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0639_ : _3488_;
  assign _3489_ = _0977_[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) datin_buf_2d[111:84] : mem_data6[111:84];
  assign _1987_[27:0] = _2668_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0647_ : _3489_;
  assign _3490_ = _0977_[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) datin_buf_2d[111:84] : mem_data7[111:84];
  assign _1988_[27:0] = _2669_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3605" *) _0655_ : _3490_;
  assign _1989_[27:0] = _2662_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0315_ : _3483_;
  assign _3491_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1989_[27:0] : 28'b0000000000000000000000000000;
  assign _1990_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1981_[27:0] : _3491_[27:0];
  assign _0976_[111:84] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0902_ : _1990_[27:0];
  assign _1991_[27:0] = _2663_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0327_ : _3484_;
  assign _1992_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1991_[27:0] : 28'b0000000000000000000000000000;
  assign _1993_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1982_[27:0] : _1992_[27:0];
  assign _0982_[111:84] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0912_ : _1993_[27:0];
  assign _1994_[27:0] = _2664_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0339_ : _3485_;
  assign _1995_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1994_[27:0] : 28'b0000000000000000000000000000;
  assign _1996_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1983_[27:0] : _1995_[27:0];
  assign _0985_[111:84] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0922_ : _1996_[27:0];
  assign _1997_[27:0] = _2665_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0351_ : _3486_;
  assign _1998_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1997_[27:0] : 28'b0000000000000000000000000000;
  assign _1999_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1984_[27:0] : _1998_[27:0];
  assign _0988_[111:84] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0932_ : _1999_[27:0];
  assign _2000_[27:0] = _2666_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0363_ : _3487_;
  assign _2001_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _2000_[27:0] : 28'b0000000000000000000000000000;
  assign _2002_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1985_[27:0] : _2001_[27:0];
  assign _0991_[111:84] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0942_ : _2002_[27:0];
  assign _2003_[27:0] = _2667_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0375_ : _3488_;
  assign _2004_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _2003_[27:0] : 28'b0000000000000000000000000000;
  assign _2005_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1986_[27:0] : _2004_[27:0];
  assign _0994_[111:84] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0952_ : _2005_[27:0];
  assign _2006_[27:0] = _2668_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0387_ : _3489_;
  assign _2007_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _2006_[27:0] : 28'b0000000000000000000000000000;
  assign _2008_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1987_[27:0] : _2007_[27:0];
  assign _0997_[111:84] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0962_ : _2008_[27:0];
  assign _2009_[27:0] = _2669_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0399_ : _3490_;
  assign _2010_[27:0] = _0979_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _2009_[27:0] : 28'b0000000000000000000000000000;
  assign _3492_[27:0] = _0980_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _1988_[27:0] : _2010_[27:0];
  assign _1000_[111:84] = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3606" *) _0972_ : _3492_[27:0];
  assign _3493_[111:0] = mem_re_1st_d[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3645" *) datin_buf : mem_rdata_0[111:0];
  assign _3494_[111:0] = mem_re_1st_d[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3646" *) datin_buf : mem_rdata_1[111:0];
  assign _3495_[111:0] = mem_re_1st_d[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3647" *) datin_buf : mem_rdata_2[111:0];
  assign _3496_[111:0] = mem_re_1st_d[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3648" *) datin_buf : mem_rdata_3[111:0];
  assign _3497_[111:0] = mem_re_1st_d[4] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3649" *) datin_buf : mem_rdata_4[111:0];
  assign _3498_[111:0] = mem_re_1st_d[5] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3650" *) datin_buf : mem_rdata_5[111:0];
  assign _3499_[111:0] = mem_re_1st_d[6] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3651" *) datin_buf : mem_rdata_6[111:0];
  assign _3500_[111:0] = mem_re_1st_d[7] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:3652" *) datin_buf : mem_rdata_7[111:0];
  assign pooling1d_vld_rebuild = _2670_ ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4333" *) 1'b1 : pooling1d_pvld;
  assign mem_data_valid = load_wr_stage2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4384" *) mem_re_2d : 8'b00000000;
  assign pooling_2d_result_0 = mem_re_1st_2d[0] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4393" *) datin_buf_2d : _0976_;
  assign pooling_2d_result_1 = mem_re_1st_2d[1] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4394" *) datin_buf_2d : _0982_;
  assign pooling_2d_result_2 = mem_re_1st_2d[2] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4395" *) datin_buf_2d : _0985_;
  assign pooling_2d_result_3 = mem_re_1st_2d[3] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4396" *) datin_buf_2d : _0988_;
  assign pooling_2d_result_4 = mem_re_1st_2d[4] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4397" *) datin_buf_2d : _0991_;
  assign pooling_2d_result_5 = mem_re_1st_2d[5] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4398" *) datin_buf_2d : _0994_;
  assign pooling_2d_result_6 = mem_re_1st_2d[6] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4399" *) datin_buf_2d : _0997_;
  assign pooling_2d_result_7 = mem_re_1st_2d[7] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4400" *) datin_buf_2d : _1000_;
  assign mem_wdata_0 = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4558" *) { din_pd_d4[132:129], 11'b00000000000, fp_mem0_wdata[100:0] } : int_mem_wdata_0;
  assign mem_wdata_1 = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4559" *) { din_pd_d4[136:133], 11'b00000000000, fp_mem1_wdata[100:0] } : int_mem_wdata_1;
  assign mem_wdata_2 = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4560" *) { din_pd_d4[140:137], 11'b00000000000, fp_mem2_wdata[100:0] } : int_mem_wdata_2;
  assign mem_wdata_3 = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4561" *) { din_pd_d4[144:141], 11'b00000000000, fp_mem3_wdata[100:0] } : int_mem_wdata_3;
  assign mem_wdata_4 = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4562" *) { din_pd_d4[148:145], 11'b00000000000, fp_mem4_wdata[100:0] } : int_mem_wdata_4;
  assign mem_wdata_5 = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4563" *) { din_pd_d4[152:149], 11'b00000000000, fp_mem5_wdata[100:0] } : int_mem_wdata_5;
  assign mem_wdata_6 = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4564" *) { din_pd_d4[156:153], 11'b00000000000, fp_mem6_wdata[100:0] } : int_mem_wdata_6;
  assign mem_wdata_7 = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4565" *) { din_pd_d4[160:157], 11'b00000000000, fp_mem7_wdata[100:0] } : int_mem_wdata_7;
  assign mem_we = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4566" *) fp_mem_we : _1709_;
  assign mem_waddr_0 = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4567" *) din_pd_d4[120:115] : int_mem_waddr;
  assign wr_data_stage1_prdy = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:5847" *) fp16_add_in_rdy : _2693_;
  assign pout_mem_data = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6193" *) fp16_mul_pad_line_in_pd_d3 : int_pout_mem_data;
  assign pout_mem_size_v_use = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6219" *) fp16_mul_pad_line_in_pd_d0[114:112] : pout_mem_size_v;
  assign data_16bit_0 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6298" *) data_16bit_0_ff : pout_mem_data_0[21:0];
  assign data_16bit_1 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6299" *) data_16bit_1_ff : pout_mem_data_1[21:0];
  assign data_16bit_2 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6300" *) data_16bit_2_ff : pout_mem_data_2[21:0];
  assign data_16bit_3 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6301" *) data_16bit_3_ff : pout_mem_data_3[21:0];
  assign data_8bit_0 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6310" *) data_8bit_0_ff : pout_mem_data_0[13:0];
  assign data_8bit_1 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6311" *) data_8bit_1_ff : pout_mem_data_0[27:14];
  assign data_8bit_2 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6312" *) data_8bit_2_ff : pout_mem_data_1[13:0];
  assign data_8bit_3 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6313" *) data_8bit_3_ff : pout_mem_data_1[27:14];
  assign data_8bit_4 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6314" *) data_8bit_4_ff : pout_mem_data_2[13:0];
  assign data_8bit_5 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6315" *) data_8bit_5_ff : pout_mem_data_2[27:14];
  assign data_8bit_6 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6316" *) data_8bit_6_ff : pout_mem_data_3[13:0];
  assign data_8bit_7 = padding_here ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6317" *) data_8bit_7_ff : pout_mem_data_3[27:14];
  assign data_hmult_16bit_0_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6370" *) data_hmult_16bit_0_ext_ff : { pout_data_0_0[21], pout_data_0_0[21:0], 16'b0000000000000000 };
  assign data_hmult_16bit_1_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6371" *) data_hmult_16bit_1_ext_ff : { pout_data_0_1[21], pout_data_0_1[21:0], 16'b0000000000000000 };
  assign data_hmult_16bit_2_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6372" *) data_hmult_16bit_2_ext_ff : { pout_data_0_2[21], pout_data_0_2[21:0], 16'b0000000000000000 };
  assign data_hmult_16bit_3_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6373" *) data_hmult_16bit_3_ext_ff : { pout_data_0_3[21], pout_data_0_3[21:0], 16'b0000000000000000 };
  assign _3501_ = i16_more_neg_0_5_0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6386" *) i16_neg_add1_0 : _1265_;
  assign data_hmult_16bit_0 = i16_less_neg_0_5_0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6386" *) data_hmult_16bit_0_ext[34:16] : _3501_;
  assign _3502_ = i16_more_neg_0_5_1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6387" *) i16_neg_add1_1 : _1266_;
  assign data_hmult_16bit_1 = i16_less_neg_0_5_1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6387" *) data_hmult_16bit_1_ext[34:16] : _3502_;
  assign _3503_ = i16_more_neg_0_5_2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6388" *) i16_neg_add1_2 : _1267_;
  assign data_hmult_16bit_2 = i16_less_neg_0_5_2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6388" *) data_hmult_16bit_2_ext[34:16] : _3503_;
  assign _3504_ = i16_more_neg_0_5_3 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6389" *) i16_neg_add1_3 : _1268_;
  assign data_hmult_16bit_3 = i16_less_neg_0_5_3 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6389" *) data_hmult_16bit_3_ext[34:16] : _3504_;
  assign data_hmult_8bit_0_lsb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6579" *) data_hmult_8bit_0_lsb_ext_ff : { pout_data_0_0[13], pout_data_0_0[13:0], 16'b0000000000000000 };
  assign data_hmult_8bit_0_msb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6580" *) data_hmult_8bit_0_msb_ext_ff : { pout_data_0_0[27], pout_data_0_0[27:14], 16'b0000000000000000 };
  assign data_hmult_8bit_1_lsb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6581" *) data_hmult_8bit_1_lsb_ext_ff : { pout_data_0_1[13], pout_data_0_1[13:0], 16'b0000000000000000 };
  assign data_hmult_8bit_1_msb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6582" *) data_hmult_8bit_1_msb_ext_ff : { pout_data_0_1[27], pout_data_0_1[27:14], 16'b0000000000000000 };
  assign data_hmult_8bit_2_lsb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6583" *) data_hmult_8bit_2_lsb_ext_ff : { pout_data_0_2[13], pout_data_0_2[13:0], 16'b0000000000000000 };
  assign data_hmult_8bit_2_msb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6584" *) data_hmult_8bit_2_msb_ext_ff : { pout_data_0_2[27], pout_data_0_2[27:14], 16'b0000000000000000 };
  assign data_hmult_8bit_3_lsb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6585" *) data_hmult_8bit_3_lsb_ext_ff : { pout_data_0_3[13], pout_data_0_3[13:0], 16'b0000000000000000 };
  assign data_hmult_8bit_3_msb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6586" *) data_hmult_8bit_3_msb_ext_ff : { pout_data_0_3[27], pout_data_0_3[27:14], 16'b0000000000000000 };
  assign _3505_ = i8_more_neg_0_5_0_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6611" *) i8_neg_add1_0_l : _1269_;
  assign hmult_8bit_0_lsb = i8_less_neg_0_5_0_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6611" *) data_hmult_8bit_0_lsb_ext[26:16] : _3505_;
  assign _3506_ = i8_more_neg_0_5_0_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6612" *) i8_neg_add1_0_m : _1270_;
  assign hmult_8bit_0_msb = i8_less_neg_0_5_0_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6612" *) data_hmult_8bit_0_msb_ext[26:16] : _3506_;
  assign _3507_ = i8_more_neg_0_5_1_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6613" *) i8_neg_add1_1_l : _1271_;
  assign hmult_8bit_1_lsb = i8_less_neg_0_5_1_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6613" *) data_hmult_8bit_1_lsb_ext[26:16] : _3507_;
  assign _3508_ = i8_more_neg_0_5_1_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6614" *) i8_neg_add1_1_m : _1272_;
  assign hmult_8bit_1_msb = i8_less_neg_0_5_1_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6614" *) data_hmult_8bit_1_msb_ext[26:16] : _3508_;
  assign _3509_ = i8_more_neg_0_5_2_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6615" *) i8_neg_add1_2_l : _1273_;
  assign hmult_8bit_2_lsb = i8_less_neg_0_5_2_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6615" *) data_hmult_8bit_2_lsb_ext[26:16] : _3509_;
  assign _3510_ = i8_more_neg_0_5_2_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6616" *) i8_neg_add1_2_m : _1274_;
  assign hmult_8bit_2_msb = i8_less_neg_0_5_2_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6616" *) data_hmult_8bit_2_msb_ext[26:16] : _3510_;
  assign _3511_ = i8_more_neg_0_5_3_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6617" *) i8_neg_add1_3_l : _1275_;
  assign hmult_8bit_3_lsb = i8_less_neg_0_5_3_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6617" *) data_hmult_8bit_3_lsb_ext[26:16] : _3511_;
  assign _3512_ = i8_more_neg_0_5_3_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6618" *) i8_neg_add1_3_m : _1276_;
  assign hmult_8bit_3_msb = i8_less_neg_0_5_3_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6618" *) data_hmult_8bit_3_msb_ext[26:16] : _3512_;
  assign data_hmult_stage0_in0 = int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6983" *) { hmult_8bit_0_msb, hmult_8bit_0_lsb } : { data_hmult_16bit_0[18], data_hmult_16bit_0[18], data_hmult_16bit_0[18], data_hmult_16bit_0 };
  assign data_hmult_stage0_in1 = int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6984" *) { hmult_8bit_1_msb, hmult_8bit_1_lsb } : { data_hmult_16bit_1[18], data_hmult_16bit_1[18], data_hmult_16bit_1[18], data_hmult_16bit_1 };
  assign data_hmult_stage0_in2 = int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6985" *) { hmult_8bit_2_msb, hmult_8bit_2_lsb } : { data_hmult_16bit_2[18], data_hmult_16bit_2[18], data_hmult_16bit_2[18], data_hmult_16bit_2 };
  assign data_hmult_stage0_in3 = int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:6986" *) { hmult_8bit_3_msb, hmult_8bit_3_lsb } : { data_hmult_16bit_3[18], data_hmult_16bit_3[18], data_hmult_16bit_3[18], data_hmult_16bit_3 };
  assign data_vmult_16bit_0_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7025" *) data_vmult_16bit_0_ext_ff : { pout_data_stage0_0[18], pout_data_stage0_0[18:0], 16'b0000000000000000 };
  assign data_vmult_16bit_1_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7026" *) data_vmult_16bit_1_ext_ff : { pout_data_stage0_1[18], pout_data_stage0_1[18:0], 16'b0000000000000000 };
  assign data_vmult_16bit_2_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7027" *) data_vmult_16bit_2_ext_ff : { pout_data_stage0_2[18], pout_data_stage0_2[18:0], 16'b0000000000000000 };
  assign data_vmult_16bit_3_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7028" *) data_vmult_16bit_3_ext_ff : { pout_data_stage0_3[18], pout_data_stage0_3[18:0], 16'b0000000000000000 };
  assign _3513_ = i16_vmore_neg_0_5_0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7041" *) i16_neg_vadd1_0 : _1277_;
  assign data_vmult_16bit_0 = i16_vless_neg_0_5_0 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7041" *) data_vmult_16bit_0_ext[31:16] : _3513_;
  assign _3514_ = i16_vmore_neg_0_5_1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7042" *) i16_neg_vadd1_1 : _1278_;
  assign data_vmult_16bit_1 = i16_vless_neg_0_5_1 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7042" *) data_vmult_16bit_1_ext[31:16] : _3514_;
  assign _3515_ = i16_vmore_neg_0_5_2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7043" *) i16_neg_vadd1_2 : _1279_;
  assign data_vmult_16bit_2 = i16_vless_neg_0_5_2 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7043" *) data_vmult_16bit_2_ext[31:16] : _3515_;
  assign _3516_ = i16_vmore_neg_0_5_3 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7044" *) i16_neg_vadd1_3 : _1280_;
  assign data_vmult_16bit_3 = i16_vless_neg_0_5_3 ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7044" *) data_vmult_16bit_3_ext[31:16] : _3516_;
  assign data_vmult_8bit_0_lsb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7234" *) data_vmult_8bit_0_lsb_ext_ff : { pout_data_stage0_0[10], pout_data_stage0_0[10:0], 16'b0000000000000000 };
  assign data_vmult_8bit_0_msb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7235" *) data_vmult_8bit_0_msb_ext_ff : { pout_data_stage0_0[21], pout_data_stage0_0[21:11], 16'b0000000000000000 };
  assign data_vmult_8bit_1_lsb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7236" *) data_vmult_8bit_1_lsb_ext_ff : { pout_data_stage0_1[10], pout_data_stage0_1[10:0], 16'b0000000000000000 };
  assign data_vmult_8bit_1_msb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7237" *) data_vmult_8bit_1_msb_ext_ff : { pout_data_stage0_1[21], pout_data_stage0_1[21:11], 16'b0000000000000000 };
  assign data_vmult_8bit_2_lsb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7238" *) data_vmult_8bit_2_lsb_ext_ff : { pout_data_stage0_2[10], pout_data_stage0_2[10:0], 16'b0000000000000000 };
  assign data_vmult_8bit_2_msb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7239" *) data_vmult_8bit_2_msb_ext_ff : { pout_data_stage0_2[21], pout_data_stage0_2[21:11], 16'b0000000000000000 };
  assign data_vmult_8bit_3_lsb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7240" *) data_vmult_8bit_3_lsb_ext_ff : { pout_data_stage0_3[10], pout_data_stage0_3[10:0], 16'b0000000000000000 };
  assign data_vmult_8bit_3_msb_ext = average_pooling_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7241" *) data_vmult_8bit_3_msb_ext_ff : { pout_data_stage0_3[21], pout_data_stage0_3[21:11], 16'b0000000000000000 };
  assign _3517_ = i8_vmore_neg_0_5_0_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7266" *) i8_neg_vadd1_0_l : _1281_;
  assign vmult_8bit_0_lsb = i8_vless_neg_0_5_0_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7266" *) data_vmult_8bit_0_lsb_ext[23:16] : _3517_;
  assign _3518_ = i8_vmore_neg_0_5_0_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7267" *) i8_neg_vadd1_0_m : _1282_;
  assign vmult_8bit_0_msb = i8_vless_neg_0_5_0_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7267" *) data_vmult_8bit_0_msb_ext[23:16] : _3518_;
  assign _3519_ = i8_vmore_neg_0_5_1_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7268" *) i8_neg_vadd1_1_l : _1283_;
  assign vmult_8bit_1_lsb = i8_vless_neg_0_5_1_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7268" *) data_vmult_8bit_1_lsb_ext[23:16] : _3519_;
  assign _3520_ = i8_vmore_neg_0_5_1_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7269" *) i8_neg_vadd1_1_m : _1284_;
  assign vmult_8bit_1_msb = i8_vless_neg_0_5_1_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7269" *) data_vmult_8bit_1_msb_ext[23:16] : _3520_;
  assign _3521_ = i8_vmore_neg_0_5_2_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7270" *) i8_neg_vadd1_2_l : _1285_;
  assign vmult_8bit_2_lsb = i8_vless_neg_0_5_2_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7270" *) data_vmult_8bit_2_lsb_ext[23:16] : _3521_;
  assign _3522_ = i8_vmore_neg_0_5_2_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7271" *) i8_neg_vadd1_2_m : _1286_;
  assign vmult_8bit_2_msb = i8_vless_neg_0_5_2_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7271" *) data_vmult_8bit_2_msb_ext[23:16] : _3522_;
  assign _3523_ = i8_vmore_neg_0_5_3_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7272" *) i8_neg_vadd1_3_l : _1287_;
  assign vmult_8bit_3_lsb = i8_vless_neg_0_5_3_l ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7272" *) data_vmult_8bit_3_lsb_ext[23:16] : _3523_;
  assign _3524_ = i8_vmore_neg_0_5_3_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7273" *) i8_neg_vadd1_3_m : _1288_;
  assign vmult_8bit_3_msb = i8_vless_neg_0_5_3_m ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7273" *) data_vmult_8bit_3_msb_ext[23:16] : _3524_;
  assign data_mult_stage1_in0 = int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7638" *) { vmult_8bit_0_msb, vmult_8bit_0_lsb } : data_vmult_16bit_0;
  assign data_mult_stage1_in1 = int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7639" *) { vmult_8bit_1_msb, vmult_8bit_1_lsb } : data_vmult_16bit_1;
  assign data_mult_stage1_in2 = int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7640" *) { vmult_8bit_2_msb, vmult_8bit_2_lsb } : data_vmult_16bit_2;
  assign data_mult_stage1_in3 = int8_en ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7641" *) { vmult_8bit_3_msb, vmult_8bit_3_lsb } : data_vmult_16bit_3;
  assign pout_data_stage3_prdy = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7675" *) 1'b0 : pdp_dp2wdma_ready;
  assign fp_mem0_wdata[100:0] = din_pd_d4[169] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7967" *) { din_pd_d4[244:228], 11'b00000000000, din_pd_d4[227:211], 11'b00000000000, din_pd_d4[210:194], 11'b00000000000, din_pd_d4[193:177] } : { fp_pooling_result_dp_0[67:51], 11'b00000000000, fp_pooling_result_dp_0[50:34], 11'b00000000000, fp_pooling_result_dp_0[33:17], 11'b00000000000, fp_pooling_result_dp_0[16:0] };
  assign fp_mem1_wdata[100:0] = din_pd_d4[170] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7972" *) { din_pd_d4[244:228], 11'b00000000000, din_pd_d4[227:211], 11'b00000000000, din_pd_d4[210:194], 11'b00000000000, din_pd_d4[193:177] } : { fp_pooling_result_dp_1[67:51], 11'b00000000000, fp_pooling_result_dp_1[50:34], 11'b00000000000, fp_pooling_result_dp_1[33:17], 11'b00000000000, fp_pooling_result_dp_1[16:0] };
  assign fp_mem2_wdata[100:0] = din_pd_d4[171] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7977" *) { din_pd_d4[244:228], 11'b00000000000, din_pd_d4[227:211], 11'b00000000000, din_pd_d4[210:194], 11'b00000000000, din_pd_d4[193:177] } : { fp_pooling_result_dp_2[67:51], 11'b00000000000, fp_pooling_result_dp_2[50:34], 11'b00000000000, fp_pooling_result_dp_2[33:17], 11'b00000000000, fp_pooling_result_dp_2[16:0] };
  assign fp_mem3_wdata[100:0] = din_pd_d4[172] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7982" *) { din_pd_d4[244:228], 11'b00000000000, din_pd_d4[227:211], 11'b00000000000, din_pd_d4[210:194], 11'b00000000000, din_pd_d4[193:177] } : { fp_pooling_result_dp_3[67:51], 11'b00000000000, fp_pooling_result_dp_3[50:34], 11'b00000000000, fp_pooling_result_dp_3[33:17], 11'b00000000000, fp_pooling_result_dp_3[16:0] };
  assign fp_mem4_wdata[100:0] = din_pd_d4[173] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7987" *) { din_pd_d4[244:228], 11'b00000000000, din_pd_d4[227:211], 11'b00000000000, din_pd_d4[210:194], 11'b00000000000, din_pd_d4[193:177] } : { fp_pooling_result_dp_4[67:51], 11'b00000000000, fp_pooling_result_dp_4[50:34], 11'b00000000000, fp_pooling_result_dp_4[33:17], 11'b00000000000, fp_pooling_result_dp_4[16:0] };
  assign fp_mem5_wdata[100:0] = din_pd_d4[174] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7992" *) { din_pd_d4[244:228], 11'b00000000000, din_pd_d4[227:211], 11'b00000000000, din_pd_d4[210:194], 11'b00000000000, din_pd_d4[193:177] } : { fp_pooling_result_dp_5[67:51], 11'b00000000000, fp_pooling_result_dp_5[50:34], 11'b00000000000, fp_pooling_result_dp_5[33:17], 11'b00000000000, fp_pooling_result_dp_5[16:0] };
  assign fp_mem6_wdata[100:0] = din_pd_d4[175] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7997" *) { din_pd_d4[244:228], 11'b00000000000, din_pd_d4[227:211], 11'b00000000000, din_pd_d4[210:194], 11'b00000000000, din_pd_d4[193:177] } : { fp_pooling_result_dp_6[67:51], 11'b00000000000, fp_pooling_result_dp_6[50:34], 11'b00000000000, fp_pooling_result_dp_6[33:17], 11'b00000000000, fp_pooling_result_dp_6[16:0] };
  assign fp_mem7_wdata[100:0] = din_pd_d4[176] ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8002" *) { din_pd_d4[244:228], 11'b00000000000, din_pd_d4[227:211], 11'b00000000000, din_pd_d4[210:194], 11'b00000000000, din_pd_d4[193:177] } : { fp_pooling_result_dp_7[67:51], 11'b00000000000, fp_pooling_result_dp_7[50:34], 11'b00000000000, fp_pooling_result_dp_7[33:17], 11'b00000000000, fp_pooling_result_dp_7[16:0] };
  assign _3525_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8023" *) _1895_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3526_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8024" *) _1896_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3527_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8025" *) _1897_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3528_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8026" *) _1898_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3529_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8027" *) _1899_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3530_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8028" *) _1900_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3531_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8029" *) _1901_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3532_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8030" *) _1902_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3533_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8031" *) _1903_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3534_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8032" *) _1904_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3535_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8033" *) _1905_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3536_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8034" *) _1906_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3537_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8035" *) _1907_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3538_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8036" *) _1908_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3539_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8037" *) _1909_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _3540_ = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8038" *) _1910_ : 115'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign fp16_mulw_in_vld = fp_add_out_vld ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8762" *) _3138_ : 1'b0;
  assign pdp_dp2wdma_pd = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9111" *) { fp17T16_out3, fp17T16_out2, fp17T16_out1, fp17T16_out0 } : { pout_data_stage1_3, pout_data_stage1_2, pout_data_stage1_1, pout_data_stage1_0 };
  assign pdp_dp2wdma_valid = fp16_mean_pool_cfg ? (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9112" *) fp_dp2wdma_pvld : int_dp2wdma_valid;
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4579" *)
  nv_ram_rws_64x116 bank0_uram_0 (
    .clk(nvdla_core_clk),
    .di(mem_wdata_0),
    .dout(mem_rdata_0),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sub_lbuf_dout_cnt),
    .re(_2671_),
    .wa(mem_waddr_0),
    .we(mem_we[0])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4589" *)
  nv_ram_rws_64x116 bank1_uram_0 (
    .clk(nvdla_core_clk),
    .di(mem_wdata_1),
    .dout(mem_rdata_1),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sub_lbuf_dout_cnt),
    .re(_2672_),
    .wa(mem_waddr_0),
    .we(mem_we[1])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4599" *)
  nv_ram_rws_64x116 bank2_uram_0 (
    .clk(nvdla_core_clk),
    .di(mem_wdata_2),
    .dout(mem_rdata_2),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sub_lbuf_dout_cnt),
    .re(_2673_),
    .wa(mem_waddr_0),
    .we(mem_we[2])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4609" *)
  nv_ram_rws_64x116 bank3_uram_0 (
    .clk(nvdla_core_clk),
    .di(mem_wdata_3),
    .dout(mem_rdata_3),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sub_lbuf_dout_cnt),
    .re(_2674_),
    .wa(mem_waddr_0),
    .we(mem_we[3])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4619" *)
  nv_ram_rws_64x116 bank4_uram_0 (
    .clk(nvdla_core_clk),
    .di(mem_wdata_4),
    .dout(mem_rdata_4),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sub_lbuf_dout_cnt),
    .re(_2675_),
    .wa(mem_waddr_0),
    .we(mem_we[4])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4629" *)
  nv_ram_rws_64x116 bank5_uram_0 (
    .clk(nvdla_core_clk),
    .di(mem_wdata_5),
    .dout(mem_rdata_5),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sub_lbuf_dout_cnt),
    .re(_2676_),
    .wa(mem_waddr_0),
    .we(mem_we[5])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4639" *)
  nv_ram_rws_64x116 bank6_uram_0 (
    .clk(nvdla_core_clk),
    .di(mem_wdata_6),
    .dout(mem_rdata_6),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sub_lbuf_dout_cnt),
    .re(_2677_),
    .wa(mem_waddr_0),
    .we(mem_we[6])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:4649" *)
  nv_ram_rws_64x116 bank7_uram_0 (
    .clk(nvdla_core_clk),
    .di(mem_wdata_7),
    .dout(mem_rdata_7),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sub_lbuf_dout_cnt),
    .re(_2678_),
    .wa(mem_waddr_0),
    .we(mem_we[7])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8793" *)
  HLS_fp17_mul mul_padx_kwidth (
    .chn_a_rsc_lz(fp16_mul_pad_line_rdy[0]),
    .chn_a_rsc_vz(fp16_mul_pad_line_vld[0]),
    .chn_a_rsc_z(pad_table_out[16:0]),
    .chn_b_rsc_lz(fp16_mul_pad_line_rdy[1]),
    .chn_b_rsc_vz(fp16_mul_pad_line_vld[1]),
    .chn_b_rsc_z(kernel_width_fp17),
    .chn_o_rsc_lz(pad_line_sum_pvld),
    .chn_o_rsc_vz(pad_line_sum_prdy),
    .chn_o_rsc_z(pad_line_sum),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7899" *)
  NV_NVDLA_PDP_CORE_CAL2D_pipe_p1 pipe_p1 (
    .din_pd_d0({ one_width_disable_2d, mem_re_2d, cur_datin_disable_2d, datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0], mem_re_1st_2d, pout_mem_data_sel_last, wr_line_end_2d, mem_data7[114:112], wr_line_end_2d, mem_data6[114:112], wr_line_end_2d, mem_data5[114:112], wr_line_end_2d, mem_data4[114:112], wr_line_end_2d, mem_data3[114:112], wr_line_end_2d, mem_data2[114:112], wr_line_end_2d, mem_data1[114:112], wr_line_end_2d, mem_data0[114:112], pout_mem_data_sel, mem_raddr_2d, pout_mem_data_last }),
    .din_pd_d1(din_pd_d1),
    .din_rdy_d0(din_rdy),
    .din_rdy_d1(din_rdy_d1),
    .din_vld_d0(din_vld_d0),
    .din_vld_d1(din_vld_d1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .nvdla_op_gated_clk_fp16(nvdla_op_gated_clk_fp16)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7909" *)
  NV_NVDLA_PDP_CORE_CAL2D_pipe_p2 pipe_p2 (
    .din_pd_d1(din_pd_d1),
    .din_pd_d2(din_pd_d2),
    .din_rdy_d1(din_rdy_d1),
    .din_rdy_d2(din_rdy_d2),
    .din_vld_d1(din_vld_d1),
    .din_vld_d2(din_vld_d2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .nvdla_op_gated_clk_fp16(nvdla_op_gated_clk_fp16)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7919" *)
  NV_NVDLA_PDP_CORE_CAL2D_pipe_p3 pipe_p3 (
    .din_pd_d2(din_pd_d2),
    .din_pd_d3(din_pd_d3),
    .din_rdy_d2(din_rdy_d2),
    .din_rdy_d3(din_rdy_d3),
    .din_vld_d2(din_vld_d2),
    .din_vld_d3(din_vld_d3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .nvdla_op_gated_clk_fp16(nvdla_op_gated_clk_fp16)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7929" *)
  NV_NVDLA_PDP_CORE_CAL2D_pipe_p4 pipe_p4 (
    .din_pd_d3(din_pd_d3),
    .din_pd_d4(din_pd_d4),
    .din_rdy_d3(din_rdy_d3),
    .din_rdy_d4(din_rdy_d4),
    .din_vld_d3(din_vld_d3),
    .din_vld_d4(din_vld_d4),
    .nvdla_core_rstn(nvdla_core_rstn),
    .nvdla_op_gated_clk_fp16(nvdla_op_gated_clk_fp16)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8809" *)
  NV_NVDLA_PDP_CORE_CAL2D_pipe_p5 pipe_p5 (
    .fp16_mul_pad_line_in_pd_d0(fp16_mul_pad_line_in_pd_d0),
    .fp16_mul_pad_line_in_pd_d1(fp16_mul_pad_line_in_pd_d1),
    .fp16_mul_pad_line_in_rdy_d0(fp16_mul_pad_line_in_rdy),
    .fp16_mul_pad_line_in_rdy_d1(fp16_mul_pad_line_in_rdy_d1),
    .fp16_mul_pad_line_in_vld_d0(fp16_mul_pad_line_in_vld_d0),
    .fp16_mul_pad_line_in_vld_d1(fp16_mul_pad_line_in_vld_d1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .nvdla_op_gated_clk_fp16(nvdla_op_gated_clk_fp16)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8819" *)
  NV_NVDLA_PDP_CORE_CAL2D_pipe_p6 pipe_p6 (
    .fp16_mul_pad_line_in_pd_d1(fp16_mul_pad_line_in_pd_d1),
    .fp16_mul_pad_line_in_pd_d2(fp16_mul_pad_line_in_pd_d2),
    .fp16_mul_pad_line_in_rdy_d1(fp16_mul_pad_line_in_rdy_d1),
    .fp16_mul_pad_line_in_rdy_d2(fp16_mul_pad_line_in_rdy_d2),
    .fp16_mul_pad_line_in_vld_d1(fp16_mul_pad_line_in_vld_d1),
    .fp16_mul_pad_line_in_vld_d2(fp16_mul_pad_line_in_vld_d2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .nvdla_op_gated_clk_fp16(nvdla_op_gated_clk_fp16)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8829" *)
  NV_NVDLA_PDP_CORE_CAL2D_pipe_p7 pipe_p7 (
    .fp16_mul_pad_line_in_pd_d2(fp16_mul_pad_line_in_pd_d2),
    .fp16_mul_pad_line_in_pd_d3(fp16_mul_pad_line_in_pd_d3),
    .fp16_mul_pad_line_in_rdy_d2(fp16_mul_pad_line_in_rdy_d2),
    .fp16_mul_pad_line_in_rdy_d3(fp16_mul_pad_line_in_rdy_d3),
    .fp16_mul_pad_line_in_vld_d2(fp16_mul_pad_line_in_vld_d2),
    .fp16_mul_pad_line_in_vld_d3(fp16_mul_pad_line_in_vld_d3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .nvdla_op_gated_clk_fp16(nvdla_op_gated_clk_fp16)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8858" *)
  HLS_fp17_add u_HLS_fp17_add_0 (
    .chn_a_rsc_lz(fp16_add_pad_in_a_rdy[0]),
    .chn_a_rsc_vz(fp16_add_pad_in_a_vld[0]),
    .chn_a_rsc_z(fp16_mul_pad_line_in_pd_d3[16:0]),
    .chn_b_rsc_lz(fp16_add_pad_in_b_rdy[0]),
    .chn_b_rsc_vz(fp16_add_pad_in_b_vld[0]),
    .chn_b_rsc_z(pad_line_sum),
    .chn_o_rsc_lz(fp16_add_pad_out_vld[0]),
    .chn_o_rsc_vz(fp16_add_pad_out_rdy[0]),
    .chn_o_rsc_z(fp16_add_pad_out0),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8871" *)
  HLS_fp17_add u_HLS_fp17_add_1 (
    .chn_a_rsc_lz(fp16_add_pad_in_a_rdy[1]),
    .chn_a_rsc_vz(fp16_add_pad_in_a_vld[1]),
    .chn_a_rsc_z(fp16_mul_pad_line_in_pd_d3[44:28]),
    .chn_b_rsc_lz(fp16_add_pad_in_b_rdy[1]),
    .chn_b_rsc_vz(fp16_add_pad_in_b_vld[1]),
    .chn_b_rsc_z(pad_line_sum),
    .chn_o_rsc_lz(fp16_add_pad_out_vld[1]),
    .chn_o_rsc_vz(fp16_add_pad_out_rdy[1]),
    .chn_o_rsc_z(fp16_add_pad_out1),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8884" *)
  HLS_fp17_add u_HLS_fp17_add_2 (
    .chn_a_rsc_lz(fp16_add_pad_in_a_rdy[2]),
    .chn_a_rsc_vz(fp16_add_pad_in_a_vld[2]),
    .chn_a_rsc_z(fp16_mul_pad_line_in_pd_d3[72:56]),
    .chn_b_rsc_lz(fp16_add_pad_in_b_rdy[2]),
    .chn_b_rsc_vz(fp16_add_pad_in_b_vld[2]),
    .chn_b_rsc_z(pad_line_sum),
    .chn_o_rsc_lz(fp16_add_pad_out_vld[2]),
    .chn_o_rsc_vz(fp16_add_pad_out_rdy[2]),
    .chn_o_rsc_z(fp16_add_pad_out2),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8897" *)
  HLS_fp17_add u_HLS_fp17_add_3 (
    .chn_a_rsc_lz(fp16_add_pad_in_a_rdy[3]),
    .chn_a_rsc_vz(fp16_add_pad_in_a_vld[3]),
    .chn_a_rsc_z(fp16_mul_pad_line_in_pd_d3[100:84]),
    .chn_b_rsc_lz(fp16_add_pad_in_b_rdy[3]),
    .chn_b_rsc_vz(fp16_add_pad_in_b_vld[3]),
    .chn_b_rsc_z(pad_line_sum),
    .chn_o_rsc_lz(fp16_add_pad_out_vld[3]),
    .chn_o_rsc_vz(fp16_add_pad_out_rdy[3]),
    .chn_o_rsc_z(fp16_add_pad_out3),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9003" *)
  HLS_fp17_mul u_HLS_fp17_mulv_0 (
    .chn_a_rsc_lz(fp16_mulv_in_a_rdy[0]),
    .chn_a_rsc_vz(fp16_mulv_in_a_vld[0]),
    .chn_a_rsc_z(fp16_mulw_out0),
    .chn_b_rsc_lz(fp16_mulv_in_b_rdy[0]),
    .chn_b_rsc_vz(fp16_mulv_in_b_vld[0]),
    .chn_b_rsc_z(reg2dp_recip_height_cfg),
    .chn_o_rsc_lz(fp16_mulv_out_vld[0]),
    .chn_o_rsc_vz(fp16_mulv_out_rdy[0]),
    .chn_o_rsc_z(fp16_mulv_out0),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9016" *)
  HLS_fp17_mul u_HLS_fp17_mulv_1 (
    .chn_a_rsc_lz(fp16_mulv_in_a_rdy[1]),
    .chn_a_rsc_vz(fp16_mulv_in_a_vld[1]),
    .chn_a_rsc_z(fp16_mulw_out1),
    .chn_b_rsc_lz(fp16_mulv_in_b_rdy[1]),
    .chn_b_rsc_vz(fp16_mulv_in_b_vld[1]),
    .chn_b_rsc_z(reg2dp_recip_height_cfg),
    .chn_o_rsc_lz(fp16_mulv_out_vld[1]),
    .chn_o_rsc_vz(fp16_mulv_out_rdy[1]),
    .chn_o_rsc_z(fp16_mulv_out1),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9029" *)
  HLS_fp17_mul u_HLS_fp17_mulv_2 (
    .chn_a_rsc_lz(fp16_mulv_in_a_rdy[2]),
    .chn_a_rsc_vz(fp16_mulv_in_a_vld[2]),
    .chn_a_rsc_z(fp16_mulw_out2),
    .chn_b_rsc_lz(fp16_mulv_in_b_rdy[2]),
    .chn_b_rsc_vz(fp16_mulv_in_b_vld[2]),
    .chn_b_rsc_z(reg2dp_recip_height_cfg),
    .chn_o_rsc_lz(fp16_mulv_out_vld[2]),
    .chn_o_rsc_vz(fp16_mulv_out_rdy[2]),
    .chn_o_rsc_z(fp16_mulv_out2),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9042" *)
  HLS_fp17_mul u_HLS_fp17_mulv_3 (
    .chn_a_rsc_lz(fp16_mulv_in_a_rdy[3]),
    .chn_a_rsc_vz(fp16_mulv_in_a_vld[3]),
    .chn_a_rsc_z(fp16_mulw_out3),
    .chn_b_rsc_lz(fp16_mulv_in_b_rdy[3]),
    .chn_b_rsc_vz(fp16_mulv_in_b_vld[3]),
    .chn_b_rsc_z(reg2dp_recip_height_cfg),
    .chn_o_rsc_lz(fp16_mulv_out_vld[3]),
    .chn_o_rsc_vz(fp16_mulv_out_rdy[3]),
    .chn_o_rsc_z(fp16_mulv_out3),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8931" *)
  HLS_fp17_mul u_HLS_fp17_mulw_0 (
    .chn_a_rsc_lz(fp16_mulw_in_a_rdy[0]),
    .chn_a_rsc_vz(fp16_mulw_in_a_vld[0]),
    .chn_a_rsc_z(fp16_add_pad_out0),
    .chn_b_rsc_lz(fp16_mulw_in_b_rdy[0]),
    .chn_b_rsc_vz(fp16_mulw_in_b_vld[0]),
    .chn_b_rsc_z(reg2dp_recip_width_cfg),
    .chn_o_rsc_lz(fp16_mulw_out_vld[0]),
    .chn_o_rsc_vz(fp16_mulw_out_rdy[0]),
    .chn_o_rsc_z(fp16_mulw_out0),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8944" *)
  HLS_fp17_mul u_HLS_fp17_mulw_1 (
    .chn_a_rsc_lz(fp16_mulw_in_a_rdy[1]),
    .chn_a_rsc_vz(fp16_mulw_in_a_vld[1]),
    .chn_a_rsc_z(fp16_add_pad_out1),
    .chn_b_rsc_lz(fp16_mulw_in_b_rdy[1]),
    .chn_b_rsc_vz(fp16_mulw_in_b_vld[1]),
    .chn_b_rsc_z(reg2dp_recip_width_cfg),
    .chn_o_rsc_lz(fp16_mulw_out_vld[1]),
    .chn_o_rsc_vz(fp16_mulw_out_rdy[1]),
    .chn_o_rsc_z(fp16_mulw_out1),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8957" *)
  HLS_fp17_mul u_HLS_fp17_mulw_2 (
    .chn_a_rsc_lz(fp16_mulw_in_a_rdy[2]),
    .chn_a_rsc_vz(fp16_mulw_in_a_vld[2]),
    .chn_a_rsc_z(fp16_add_pad_out2),
    .chn_b_rsc_lz(fp16_mulw_in_b_rdy[2]),
    .chn_b_rsc_vz(fp16_mulw_in_b_vld[2]),
    .chn_b_rsc_z(reg2dp_recip_width_cfg),
    .chn_o_rsc_lz(fp16_mulw_out_vld[2]),
    .chn_o_rsc_vz(fp16_mulw_out_rdy[2]),
    .chn_o_rsc_z(fp16_mulw_out2),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:8970" *)
  HLS_fp17_mul u_HLS_fp17_mulw_3 (
    .chn_a_rsc_lz(fp16_mulw_in_a_rdy[3]),
    .chn_a_rsc_vz(fp16_mulw_in_a_vld[3]),
    .chn_a_rsc_z(fp16_add_pad_out3),
    .chn_b_rsc_lz(fp16_mulw_in_b_rdy[3]),
    .chn_b_rsc_vz(fp16_mulw_in_b_vld[3]),
    .chn_b_rsc_z(reg2dp_recip_width_cfg),
    .chn_o_rsc_lz(fp16_mulw_out_vld[3]),
    .chn_o_rsc_vz(fp16_mulw_out_rdy[3]),
    .chn_o_rsc_z(fp16_mulw_out3),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9059" *)
  HLS_fp17_to_fp16 u_HLS_fp17_to_fp16_0 (
    .chn_a_rsc_lz(fp16_mulv_out_rdy[0]),
    .chn_a_rsc_vz(fp16_mulv_out_vld[0]),
    .chn_a_rsc_z(fp16_mulv_out0),
    .chn_o_rsc_lz(fp17T16_out_vld[0]),
    .chn_o_rsc_vz(fp17T16_out_rdy[0]),
    .chn_o_rsc_z(fp17T16_out0),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9069" *)
  HLS_fp17_to_fp16 u_HLS_fp17_to_fp16_1 (
    .chn_a_rsc_lz(fp16_mulv_out_rdy[1]),
    .chn_a_rsc_vz(fp16_mulv_out_vld[1]),
    .chn_a_rsc_z(fp16_mulv_out1),
    .chn_o_rsc_lz(fp17T16_out_vld[1]),
    .chn_o_rsc_vz(fp17T16_out_rdy[1]),
    .chn_o_rsc_z(fp17T16_out1),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9079" *)
  HLS_fp17_to_fp16 u_HLS_fp17_to_fp16_2 (
    .chn_a_rsc_lz(fp16_mulv_out_rdy[2]),
    .chn_a_rsc_vz(fp16_mulv_out_vld[2]),
    .chn_a_rsc_z(fp16_mulv_out2),
    .chn_o_rsc_lz(fp17T16_out_vld[2]),
    .chn_o_rsc_vz(fp17T16_out_rdy[2]),
    .chn_o_rsc_z(fp17T16_out2),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:9089" *)
  HLS_fp17_to_fp16 u_HLS_fp17_to_fp16_3 (
    .chn_a_rsc_lz(fp16_mulv_out_rdy[3]),
    .chn_a_rsc_vz(fp16_mulv_out_vld[3]),
    .chn_a_rsc_z(fp16_mulv_out3),
    .chn_o_rsc_lz(fp17T16_out_vld[3]),
    .chn_o_rsc_vz(fp17T16_out_rdy[3]),
    .chn_o_rsc_z(fp17T16_out3),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7803" *)
  fp16_4add u_fp16_cal2d_pooling_sum_0 (
    .fp16_add_in_a({ datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0] }),
    .fp16_add_in_b({ mem_data0[100:84], mem_data0[72:56], mem_data0[44:28], mem_data0[16:0] }),
    .fp16_add_in_prdy(fp16_4add_in_prdy[0]),
    .fp16_add_in_pvld(fp16_4add_in_pvld[0]),
    .fp16_add_out_dp(fp_pooling_result_dp_0),
    .fp16_add_out_prdy(fp16_4add_out_prdy[0]),
    .fp16_add_out_pvld(fp16_4add_out_pvld[0]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7814" *)
  fp16_4add u_fp16_cal2d_pooling_sum_1 (
    .fp16_add_in_a({ datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0] }),
    .fp16_add_in_b({ mem_data1[100:84], mem_data1[72:56], mem_data1[44:28], mem_data1[16:0] }),
    .fp16_add_in_prdy(fp16_4add_in_prdy[1]),
    .fp16_add_in_pvld(fp16_4add_in_pvld[1]),
    .fp16_add_out_dp(fp_pooling_result_dp_1),
    .fp16_add_out_prdy(fp16_4add_out_prdy[1]),
    .fp16_add_out_pvld(fp16_4add_out_pvld[1]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7825" *)
  fp16_4add u_fp16_cal2d_pooling_sum_2 (
    .fp16_add_in_a({ datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0] }),
    .fp16_add_in_b({ mem_data2[100:84], mem_data2[72:56], mem_data2[44:28], mem_data2[16:0] }),
    .fp16_add_in_prdy(fp16_4add_in_prdy[2]),
    .fp16_add_in_pvld(fp16_4add_in_pvld[2]),
    .fp16_add_out_dp(fp_pooling_result_dp_2),
    .fp16_add_out_prdy(fp16_4add_out_prdy[2]),
    .fp16_add_out_pvld(fp16_4add_out_pvld[2]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7836" *)
  fp16_4add u_fp16_cal2d_pooling_sum_3 (
    .fp16_add_in_a({ datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0] }),
    .fp16_add_in_b({ mem_data3[100:84], mem_data3[72:56], mem_data3[44:28], mem_data3[16:0] }),
    .fp16_add_in_prdy(fp16_4add_in_prdy[3]),
    .fp16_add_in_pvld(fp16_4add_in_pvld[3]),
    .fp16_add_out_dp(fp_pooling_result_dp_3),
    .fp16_add_out_prdy(fp16_4add_out_prdy[3]),
    .fp16_add_out_pvld(fp16_4add_out_pvld[3]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7847" *)
  fp16_4add u_fp16_cal2d_pooling_sum_4 (
    .fp16_add_in_a({ datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0] }),
    .fp16_add_in_b({ mem_data4[100:84], mem_data4[72:56], mem_data4[44:28], mem_data4[16:0] }),
    .fp16_add_in_prdy(fp16_4add_in_prdy[4]),
    .fp16_add_in_pvld(fp16_4add_in_pvld[4]),
    .fp16_add_out_dp(fp_pooling_result_dp_4),
    .fp16_add_out_prdy(fp16_4add_out_prdy[4]),
    .fp16_add_out_pvld(fp16_4add_out_pvld[4]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7858" *)
  fp16_4add u_fp16_cal2d_pooling_sum_5 (
    .fp16_add_in_a({ datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0] }),
    .fp16_add_in_b({ mem_data5[100:84], mem_data5[72:56], mem_data5[44:28], mem_data5[16:0] }),
    .fp16_add_in_prdy(fp16_4add_in_prdy[5]),
    .fp16_add_in_pvld(fp16_4add_in_pvld[5]),
    .fp16_add_out_dp(fp_pooling_result_dp_5),
    .fp16_add_out_prdy(fp16_4add_out_prdy[5]),
    .fp16_add_out_pvld(fp16_4add_out_pvld[5]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7869" *)
  fp16_4add u_fp16_cal2d_pooling_sum_6 (
    .fp16_add_in_a({ datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0] }),
    .fp16_add_in_b({ mem_data6[100:84], mem_data6[72:56], mem_data6[44:28], mem_data6[16:0] }),
    .fp16_add_in_prdy(fp16_4add_in_prdy[6]),
    .fp16_add_in_pvld(fp16_4add_in_pvld[6]),
    .fp16_add_out_dp(fp_pooling_result_dp_6),
    .fp16_add_out_prdy(fp16_4add_out_prdy[6]),
    .fp16_add_out_pvld(fp16_4add_out_pvld[6]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/pdp/NV_NVDLA_PDP_CORE_cal2d.v:7880" *)
  fp16_4add u_fp16_cal2d_pooling_sum_7 (
    .fp16_add_in_a({ datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0] }),
    .fp16_add_in_b({ mem_data7[100:84], mem_data7[72:56], mem_data7[44:28], mem_data7[16:0] }),
    .fp16_add_in_prdy(fp16_4add_in_prdy[7]),
    .fp16_add_in_pvld(fp16_4add_in_pvld[7]),
    .fp16_add_out_dp(fp_pooling_result_dp_7),
    .fp16_add_out_prdy(fp16_4add_out_prdy[7]),
    .fp16_add_out_pvld(fp16_4add_out_pvld[7]),
    .nvdla_core_clk(nvdla_op_gated_clk_fp16),
    .nvdla_core_rstn(nvdla_core_rstn)
  );
  assign _1229_[2:1] = 2'b11;
  assign _1913_[8] = 1'b0;
  assign _1914_[2:1] = 2'b00;
  assign _1915_[2] = 1'b0;
  assign _1916_[2] = 1'b0;
  assign _1917_[2:1] = 2'b00;
  assign _1918_[2] = 1'b0;
  assign _1919_[2] = 1'b0;
  assign _1920_[2:1] = 2'b00;
  assign _1921_[2] = 1'b0;
  assign _1922_[2] = 1'b0;
  assign _1923_[2:1] = 2'b00;
  assign _1924_[2] = 1'b0;
  assign _1925_[2] = 1'b0;
  assign _1926_[2:1] = 2'b00;
  assign _1927_[2] = 1'b0;
  assign _1928_[2] = 1'b0;
  assign _1929_[2:1] = 2'b00;
  assign _1930_[2] = 1'b0;
  assign _1932_[31:28] = 4'b0000;
  assign _1933_[31:28] = 4'b0000;
  assign _1934_[31:28] = 4'b0000;
  assign _1935_[31:28] = 4'b0000;
  assign _1936_[31:28] = 4'b0000;
  assign _1937_[31:28] = 4'b0000;
  assign _1938_[31:28] = 4'b0000;
  assign _1939_[31:28] = 4'b0000;
  assign _1940_[31:28] = 4'b0000;
  assign _1941_[31:28] = 4'b0000;
  assign _1942_[31:28] = 4'b0000;
  assign _1943_[31:28] = 4'b0000;
  assign _1944_[31:28] = 4'b0000;
  assign _1945_[31:28] = 4'b0000;
  assign _1946_[31:28] = 4'b0000;
  assign _1947_[31:28] = 4'b0000;
  assign _1948_[31:28] = 4'b0000;
  assign _1949_[31:28] = 4'b0000;
  assign _1950_[31:28] = 4'b0000;
  assign _1951_[31:28] = 4'b0000;
  assign _1952_[31:28] = 4'b0000;
  assign _1953_[31:28] = 4'b0000;
  assign _1954_[31:28] = 4'b0000;
  assign _1955_[31:28] = 4'b0000;
  assign _1956_[31:28] = 4'b0000;
  assign _1957_[31:28] = 4'b0000;
  assign _1958_[31:28] = 4'b0000;
  assign _1959_[31:28] = 4'b0000;
  assign _1960_[31:28] = 4'b0000;
  assign _1961_[31:28] = 4'b0000;
  assign _1962_[31:28] = 4'b0000;
  assign _1963_[31:28] = 4'b0000;
  assign _1964_[31:28] = 4'b0000;
  assign _1965_[31:28] = 4'b0000;
  assign _1966_[31:28] = 4'b0000;
  assign _1967_[31:28] = 4'b0000;
  assign _1968_[31:28] = 4'b0000;
  assign _1969_[31:28] = 4'b0000;
  assign _1970_[31:28] = 4'b0000;
  assign _1971_[31:28] = 4'b0000;
  assign _1972_[31:28] = 4'b0000;
  assign _1973_[31:28] = 4'b0000;
  assign _1974_[31:28] = 4'b0000;
  assign _1975_[31:28] = 4'b0000;
  assign _1976_[31:28] = 4'b0000;
  assign _1977_[31:28] = 4'b0000;
  assign _1978_[31:28] = 4'b0000;
  assign _1979_[31:28] = 4'b0000;
  assign _1980_[31:28] = 4'b0000;
  assign _1981_[31:28] = 4'b0000;
  assign _1982_[31:28] = 4'b0000;
  assign _1983_[31:28] = 4'b0000;
  assign _1984_[31:28] = 4'b0000;
  assign _1985_[31:28] = 4'b0000;
  assign _1986_[31:28] = 4'b0000;
  assign _1987_[31:28] = 4'b0000;
  assign _1988_[31:28] = 4'b0000;
  assign _1989_[31:28] = 4'b0000;
  assign _1990_[31:28] = 4'b0000;
  assign _1991_[31:28] = 4'b0000;
  assign _1992_[31:28] = 4'b0000;
  assign _1993_[31:28] = 4'b0000;
  assign _1994_[31:28] = 4'b0000;
  assign _1995_[31:28] = 4'b0000;
  assign _1996_[31:28] = 4'b0000;
  assign _1997_[31:28] = 4'b0000;
  assign _1998_[31:28] = 4'b0000;
  assign _1999_[31:28] = 4'b0000;
  assign _2000_[31:28] = 4'b0000;
  assign _2001_[31:28] = 4'b0000;
  assign _2002_[31:28] = 4'b0000;
  assign _2003_[31:28] = 4'b0000;
  assign _2004_[31:28] = 4'b0000;
  assign _2005_[31:28] = 4'b0000;
  assign _2006_[31:28] = 4'b0000;
  assign _2007_[31:28] = 4'b0000;
  assign _2008_[31:28] = 4'b0000;
  assign _2009_[31:28] = 4'b0000;
  assign _2010_[31:28] = 4'b0000;
  assign _3072_[9:1] = 9'b000000000;
  assign _3139_[30:10] = { _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31], _3139_[31] };
  assign _3143_[30:4] = { _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31], _3143_[31] };
  assign _3144_[30:4] = { _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31], _3144_[31] };
  assign _3145_[12:10] = 3'b000;
  assign _3146_[12:10] = 3'b000;
  assign _3420_[31:28] = 4'b0000;
  assign _3421_[31:28] = 4'b0000;
  assign _3422_[31:28] = 4'b0000;
  assign _3423_[31:28] = 4'b0000;
  assign _3424_[31:28] = 4'b0000;
  assign _3425_[31:28] = 4'b0000;
  assign _3426_[31:28] = 4'b0000;
  assign _3427_[31:28] = 4'b0000;
  assign _3428_[31:28] = 4'b0000;
  assign _3429_[31:28] = 4'b0000;
  assign _3430_[31:28] = 4'b0000;
  assign _3431_[31:28] = 4'b0000;
  assign _3432_[31:28] = 4'b0000;
  assign _3433_[31:28] = 4'b0000;
  assign _3434_[31:28] = 4'b0000;
  assign _3435_[31:28] = 4'b0000;
  assign _3444_[31:28] = 4'b0000;
  assign _3445_[31:28] = 4'b0000;
  assign _3446_[31:28] = 4'b0000;
  assign _3447_[31:28] = 4'b0000;
  assign _3448_[31:28] = 4'b0000;
  assign _3449_[31:28] = 4'b0000;
  assign _3450_[31:28] = 4'b0000;
  assign _3451_[31:28] = 4'b0000;
  assign _3452_[31:28] = 4'b0000;
  assign _3453_[31:28] = 4'b0000;
  assign _3454_[31:28] = 4'b0000;
  assign _3455_[31:28] = 4'b0000;
  assign _3456_[31:28] = 4'b0000;
  assign _3457_[31:28] = 4'b0000;
  assign _3458_[31:28] = 4'b0000;
  assign _3467_[31:28] = 4'b0000;
  assign _3468_[31:28] = 4'b0000;
  assign _3469_[31:28] = 4'b0000;
  assign _3470_[31:28] = 4'b0000;
  assign _3471_[31:28] = 4'b0000;
  assign _3472_[31:28] = 4'b0000;
  assign _3473_[31:28] = 4'b0000;
  assign _3474_[31:28] = 4'b0000;
  assign _3475_[31:28] = 4'b0000;
  assign _3476_[31:28] = 4'b0000;
  assign _3477_[31:28] = 4'b0000;
  assign _3478_[31:28] = 4'b0000;
  assign _3479_[31:28] = 4'b0000;
  assign _3480_[31:28] = 4'b0000;
  assign _3481_[31:28] = 4'b0000;
  assign _3482_[31:28] = 4'b0000;
  assign _3491_[31:28] = 4'b0000;
  assign _3492_[31:28] = 4'b0000;
  assign _3493_[114:112] = unit2d_vsize_cnt_0_d;
  assign _3494_[114:112] = unit2d_vsize_cnt_1_d;
  assign _3495_[114:112] = unit2d_vsize_cnt_2_d;
  assign _3496_[114:112] = unit2d_vsize_cnt_3_d;
  assign _3497_[114:112] = unit2d_vsize_cnt_4_d;
  assign _3498_[114:112] = unit2d_vsize_cnt_5_d;
  assign _3499_[114:112] = unit2d_vsize_cnt_6_d;
  assign _3500_[114:112] = unit2d_vsize_cnt_7_d;
  assign BANK_DEPTH = 6'b111111;
  assign buffer_lines_3 = 4'b0010;
  assign cur_datin_disable_2d_sync = din_pd_d4[245];
  assign data_hmult_8bit_0 = { hmult_8bit_0_msb, hmult_8bit_0_lsb };
  assign data_hmult_8bit_1 = { hmult_8bit_1_msb, hmult_8bit_1_lsb };
  assign data_hmult_8bit_2 = { hmult_8bit_2_msb, hmult_8bit_2_lsb };
  assign data_hmult_8bit_3 = { hmult_8bit_3_msb, hmult_8bit_3_lsb };
  assign data_vmult_8bit_0 = { vmult_8bit_0_msb, vmult_8bit_0_lsb };
  assign data_vmult_8bit_1 = { vmult_8bit_1_msb, vmult_8bit_1_lsb };
  assign data_vmult_8bit_2 = { vmult_8bit_2_msb, vmult_8bit_2_lsb };
  assign data_vmult_8bit_3 = { vmult_8bit_3_msb, vmult_8bit_3_lsb };
  assign din_pd = { one_width_disable_2d, mem_re_2d, cur_datin_disable_2d, datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0], mem_re_1st_2d, pout_mem_data_sel_last, wr_line_end_2d, mem_data7[114:112], wr_line_end_2d, mem_data6[114:112], wr_line_end_2d, mem_data5[114:112], wr_line_end_2d, mem_data4[114:112], wr_line_end_2d, mem_data3[114:112], wr_line_end_2d, mem_data2[114:112], wr_line_end_2d, mem_data1[114:112], wr_line_end_2d, mem_data0[114:112], pout_mem_data_sel, mem_raddr_2d, pout_mem_data_last };
  assign din_pd_d0 = { one_width_disable_2d, mem_re_2d, cur_datin_disable_2d, datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0], mem_re_1st_2d, pout_mem_data_sel_last, wr_line_end_2d, mem_data7[114:112], wr_line_end_2d, mem_data6[114:112], wr_line_end_2d, mem_data5[114:112], wr_line_end_2d, mem_data4[114:112], wr_line_end_2d, mem_data3[114:112], wr_line_end_2d, mem_data2[114:112], wr_line_end_2d, mem_data1[114:112], wr_line_end_2d, mem_data0[114:112], pout_mem_data_sel, mem_raddr_2d, pout_mem_data_last };
  assign din_rdy_d0 = din_rdy;
  assign din_vld = din_vld_d0;
  assign dout_pd = din_pd_d4;
  assign dout_rdy = din_rdy_d4;
  assign dout_vld = din_vld_d4;
  assign fp16_add_in_a = { datin_buf_2d[100:84], datin_buf_2d[72:56], datin_buf_2d[44:28], datin_buf_2d[16:0] };
  assign fp16_add_in_a_sync = din_pd_d4[244:177];
  assign fp16_add_in_b0 = { mem_data0[100:84], mem_data0[72:56], mem_data0[44:28], mem_data0[16:0] };
  assign fp16_add_in_b1 = { mem_data1[100:84], mem_data1[72:56], mem_data1[44:28], mem_data1[16:0] };
  assign fp16_add_in_b2 = { mem_data2[100:84], mem_data2[72:56], mem_data2[44:28], mem_data2[16:0] };
  assign fp16_add_in_b3 = { mem_data3[100:84], mem_data3[72:56], mem_data3[44:28], mem_data3[16:0] };
  assign fp16_add_in_b4 = { mem_data4[100:84], mem_data4[72:56], mem_data4[44:28], mem_data4[16:0] };
  assign fp16_add_in_b5 = { mem_data5[100:84], mem_data5[72:56], mem_data5[44:28], mem_data5[16:0] };
  assign fp16_add_in_b6 = { mem_data6[100:84], mem_data6[72:56], mem_data6[44:28], mem_data6[16:0] };
  assign fp16_add_in_b7 = { mem_data7[100:84], mem_data7[72:56], mem_data7[44:28], mem_data7[16:0] };
  assign fp16_mul_pad_line_in_pd = fp16_mul_pad_line_in_pd_d0;
  assign fp16_mul_pad_line_in_rdy_d0 = fp16_mul_pad_line_in_rdy;
  assign fp16_mul_pad_line_in_vld = fp16_mul_pad_line_in_vld_d0;
  assign fp16_mul_pad_line_out_pd = fp16_mul_pad_line_in_pd_d3;
  assign fp16_mul_pad_line_out_rdy = fp16_mul_pad_line_in_rdy_d3;
  assign fp16_mul_pad_line_out_vld = fp16_mul_pad_line_in_vld_d3;
  assign fp16_mulw_out_pvld = fp16_mulv_in_vld;
  assign fp16_pout_mem_data = fp16_mul_pad_line_in_pd_d3;
  assign fp_add_out_dp_ext_0 = { fp_pooling_result_dp_0[67:51], 11'b00000000000, fp_pooling_result_dp_0[50:34], 11'b00000000000, fp_pooling_result_dp_0[33:17], 11'b00000000000, fp_pooling_result_dp_0[16:0] };
  assign fp_add_out_dp_ext_1 = { fp_pooling_result_dp_1[67:51], 11'b00000000000, fp_pooling_result_dp_1[50:34], 11'b00000000000, fp_pooling_result_dp_1[33:17], 11'b00000000000, fp_pooling_result_dp_1[16:0] };
  assign fp_add_out_dp_ext_2 = { fp_pooling_result_dp_2[67:51], 11'b00000000000, fp_pooling_result_dp_2[50:34], 11'b00000000000, fp_pooling_result_dp_2[33:17], 11'b00000000000, fp_pooling_result_dp_2[16:0] };
  assign fp_add_out_dp_ext_3 = { fp_pooling_result_dp_3[67:51], 11'b00000000000, fp_pooling_result_dp_3[50:34], 11'b00000000000, fp_pooling_result_dp_3[33:17], 11'b00000000000, fp_pooling_result_dp_3[16:0] };
  assign fp_add_out_dp_ext_4 = { fp_pooling_result_dp_4[67:51], 11'b00000000000, fp_pooling_result_dp_4[50:34], 11'b00000000000, fp_pooling_result_dp_4[33:17], 11'b00000000000, fp_pooling_result_dp_4[16:0] };
  assign fp_add_out_dp_ext_5 = { fp_pooling_result_dp_5[67:51], 11'b00000000000, fp_pooling_result_dp_5[50:34], 11'b00000000000, fp_pooling_result_dp_5[33:17], 11'b00000000000, fp_pooling_result_dp_5[16:0] };
  assign fp_add_out_dp_ext_6 = { fp_pooling_result_dp_6[67:51], 11'b00000000000, fp_pooling_result_dp_6[50:34], 11'b00000000000, fp_pooling_result_dp_6[33:17], 11'b00000000000, fp_pooling_result_dp_6[16:0] };
  assign fp_add_out_dp_ext_7 = { fp_pooling_result_dp_7[67:51], 11'b00000000000, fp_pooling_result_dp_7[50:34], 11'b00000000000, fp_pooling_result_dp_7[33:17], 11'b00000000000, fp_pooling_result_dp_7[16:0] };
  assign fp_dp2wdma_dp = { fp17T16_out3, fp17T16_out2, fp17T16_out1, fp17T16_out0 };
  assign fp_mem0_waddr = din_pd_d4[120:115];
  assign fp_mem0_wdata[115:101] = { din_pd_d4[132:129], 11'b00000000000 };
  assign fp_mem1_waddr = din_pd_d4[120:115];
  assign fp_mem1_wdata[115:101] = { din_pd_d4[136:133], 11'b00000000000 };
  assign fp_mem2_waddr = din_pd_d4[120:115];
  assign fp_mem2_wdata[115:101] = { din_pd_d4[140:137], 11'b00000000000 };
  assign fp_mem3_waddr = din_pd_d4[120:115];
  assign fp_mem3_wdata[115:101] = { din_pd_d4[144:141], 11'b00000000000 };
  assign fp_mem4_waddr = din_pd_d4[120:115];
  assign fp_mem4_wdata[115:101] = { din_pd_d4[148:145], 11'b00000000000 };
  assign fp_mem5_waddr = din_pd_d4[120:115];
  assign fp_mem5_wdata[115:101] = { din_pd_d4[152:149], 11'b00000000000 };
  assign fp_mem6_waddr = din_pd_d4[120:115];
  assign fp_mem6_wdata[115:101] = { din_pd_d4[156:153], 11'b00000000000 };
  assign fp_mem7_waddr = din_pd_d4[120:115];
  assign fp_mem7_wdata[115:101] = { din_pd_d4[160:157], 11'b00000000000 };
  assign fp_mem_size_v = fp16_mul_pad_line_in_pd_d0[114:112];
  assign fp_pooling_result0 = { din_pd_d4[132:129], 11'b00000000000, fp_mem0_wdata[100:0] };
  assign fp_pooling_result1 = { din_pd_d4[136:133], 11'b00000000000, fp_mem1_wdata[100:0] };
  assign fp_pooling_result2 = { din_pd_d4[140:137], 11'b00000000000, fp_mem2_wdata[100:0] };
  assign fp_pooling_result3 = { din_pd_d4[144:141], 11'b00000000000, fp_mem3_wdata[100:0] };
  assign fp_pooling_result4 = { din_pd_d4[148:145], 11'b00000000000, fp_mem4_wdata[100:0] };
  assign fp_pooling_result5 = { din_pd_d4[152:149], 11'b00000000000, fp_mem5_wdata[100:0] };
  assign fp_pooling_result6 = { din_pd_d4[156:153], 11'b00000000000, fp_mem6_wdata[100:0] };
  assign fp_pooling_result7 = { din_pd_d4[160:157], 11'b00000000000, fp_mem7_wdata[100:0] };
  assign fp_pout_mem_data = fp16_mul_pad_line_in_pd_d0;
  assign fp_pout_mem_data_sel = din_pd_d4[128:121];
  assign fp_pout_mem_data_sel_last = din_pd_d4[168:161];
  assign int_dp2wdma_pd = { pout_data_stage1_3, pout_data_stage1_2, pout_data_stage1_1, pout_data_stage1_0 };
  assign mem_raddr = sub_lbuf_dout_cnt;
  assign mem_raddr_2d_sync = din_pd_d4[120:115];
  assign mem_re1_1st[6:0] = { mem_re1_1st[7], mem_re1_1st[7], mem_re1_1st[7], mem_re1_1st[7], mem_re1_1st[7], mem_re1_1st[7], mem_re1_1st[7] };
  assign { mem_re2_1st[6:4], mem_re2_1st[2:0] } = { mem_re2_1st[7], mem_re2_1st[7], mem_re2_1st[7], mem_re2_1st[3], mem_re2_1st[3], mem_re2_1st[3] };
  assign { mem_re3_1st[6], mem_re3_1st[4], mem_re3_1st[2], mem_re3_1st[0] } = { mem_re3_1st[7], mem_re3_1st[5], mem_re3_1st[3], mem_re3_1st[1] };
  assign mem_re_1st_2d_sync = din_pd_d4[176:169];
  assign mem_re_2d_sync = din_pd_d4[253:246];
  assign mem_waddr_1 = mem_waddr_0;
  assign mem_waddr_2 = mem_waddr_0;
  assign mem_waddr_3 = mem_waddr_0;
  assign mem_waddr_4 = mem_waddr_0;
  assign mem_waddr_5 = mem_waddr_0;
  assign mem_waddr_6 = mem_waddr_0;
  assign mem_waddr_7 = mem_waddr_0;
  assign mon_data_16bit_0 = 1'bx;
  assign mon_data_16bit_1 = 1'bx;
  assign mon_data_16bit_2 = 1'bx;
  assign mon_data_16bit_3 = 1'bx;
  assign mon_data_8bit_0 = 2'bxx;
  assign mon_data_8bit_0_ff[0] = mon_data_8bit_0_ff[1];
  assign mon_data_8bit_1 = 2'bxx;
  assign mon_data_8bit_1_ff[0] = mon_data_8bit_1_ff[1];
  assign mon_data_8bit_2 = 2'bxx;
  assign mon_data_8bit_2_ff[0] = mon_data_8bit_2_ff[1];
  assign mon_data_8bit_3 = 2'bxx;
  assign mon_data_8bit_3_ff[0] = mon_data_8bit_3_ff[1];
  assign mon_data_8bit_4 = 2'bxx;
  assign mon_data_8bit_4_ff[0] = mon_data_8bit_4_ff[1];
  assign mon_data_8bit_5 = 2'bxx;
  assign mon_data_8bit_5_ff[0] = mon_data_8bit_5_ff[1];
  assign mon_data_8bit_6 = 2'bxx;
  assign mon_data_8bit_6_ff[0] = mon_data_8bit_6_ff[1];
  assign mon_data_8bit_7 = 2'bxx;
  assign mon_data_8bit_7_ff[0] = mon_data_8bit_7_ff[1];
  assign mon_first_out_num = 1'bx;
  assign one_width_disable_2d_sync = din_pd_d4[254];
  assign pad_l = padding_v_cfg;
  assign pad_r = reg2dp_pad_bottom_cfg;
  assign padding_stride1_num = padding_v_cfg;
  assign padding_stride2_num = padding_v_cfg[2:1];
  assign padding_stride4_num[2:1] = 2'b00;
  assign pooling1d_pd_use = pooling1d_pd;
  assign pooling1d_prdy = pooling1d_prdy_use;
  assign pooling1d_pvld_use = pooling1d_pvld;
  assign pooling_2d_info = { wr_line_end_2d, mem_data7[114:112], wr_line_end_2d, mem_data6[114:112], wr_line_end_2d, mem_data5[114:112], wr_line_end_2d, mem_data4[114:112], wr_line_end_2d, mem_data3[114:112], wr_line_end_2d, mem_data2[114:112], wr_line_end_2d, mem_data1[114:112], wr_line_end_2d, mem_data0[114:112] };
  assign pooling_2d_info_0 = { wr_line_end_2d, mem_data0[114:112] };
  assign pooling_2d_info_1 = { wr_line_end_2d, mem_data1[114:112] };
  assign pooling_2d_info_2 = { wr_line_end_2d, mem_data2[114:112] };
  assign pooling_2d_info_3 = { wr_line_end_2d, mem_data3[114:112] };
  assign pooling_2d_info_4 = { wr_line_end_2d, mem_data4[114:112] };
  assign pooling_2d_info_5 = { wr_line_end_2d, mem_data5[114:112] };
  assign pooling_2d_info_6 = { wr_line_end_2d, mem_data6[114:112] };
  assign pooling_2d_info_7 = { wr_line_end_2d, mem_data7[114:112] };
  assign pooling_2d_info_sync = din_pd_d4[160:129];
  assign pooling_datin = datin_buf_2d;
  assign pooling_datin_ext = { din_pd_d4[244:228], 11'b00000000000, din_pd_d4[227:211], 11'b00000000000, din_pd_d4[210:194], 11'b00000000000, din_pd_d4[193:177] };
  assign pooling_size = buffer_lines_0;
  assign pooling_size_v = buffer_lines_0;
  assign pout_mem_data0 = pout_mem_data_0[21:0];
  assign pout_mem_data1 = pout_mem_data_1[21:0];
  assign pout_mem_data2 = pout_mem_data_2[21:0];
  assign pout_mem_data3 = pout_mem_data_3[21:0];
  assign pout_mem_data_last_sync = din_pd_d4[114:0];
  assign pout_mem_data_sel_last_sync = din_pd_d4[168:161];
  assign pout_mem_data_sel_sync = din_pd_d4[128:121];
  assign stride = pooling_stride_v;
  assign stride_1x = pooling_stride_v;
  assign stride_2x = { pooling_stride_v, 1'b0 };
  assign stride_4x = { pooling_stride_v, 2'b00 };
  assign unit2d_vsize1_1 = unit2d_vsize1_0;
  assign unit2d_vsize1_2 = unit2d_vsize1_0;
  assign unit2d_vsize1_3 = unit2d_vsize1_0;
  assign unit2d_vsize1_4 = unit2d_vsize1_0;
  assign unit2d_vsize1_5 = unit2d_vsize1_0;
  assign unit2d_vsize1_6 = unit2d_vsize1_0;
  assign unit2d_vsize1_7 = unit2d_vsize1_0;
  assign unit2d_vsize2_1 = unit2d_vsize2_0;
  assign unit2d_vsize2_2 = unit2d_vsize2_0;
  assign unit2d_vsize2_3 = unit2d_vsize2_0;
  assign unit2d_vsize2_5 = unit2d_vsize2_4;
  assign unit2d_vsize2_6 = unit2d_vsize2_4;
  assign unit2d_vsize2_7 = unit2d_vsize2_4;
  assign unit2d_vsize3_1 = unit2d_vsize3_0;
  assign unit2d_vsize3_3 = unit2d_vsize3_2;
  assign unit2d_vsize3_5 = unit2d_vsize3_4;
  assign unit2d_vsize3_7 = unit2d_vsize3_6;
  assign up_pnum0 = 3'b000;
endmodule
