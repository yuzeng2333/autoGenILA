module CDP_ICVT_chn_data_out_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_cdp_icvt.v:230" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_cdp_icvt.v:231" *)
  output outsig;
  assign outsig = in_0;
endmodule
