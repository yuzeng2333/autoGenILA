module FP32_TO_FP17_chn_o_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp32_to_fp17.v:155" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp32_to_fp17.v:156" *)
  output outsig;
  assign outsig = in_0;
endmodule
