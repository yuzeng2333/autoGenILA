module CSC_chn_data_out_rsci_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:496" *)
  input in_0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:497" *)
  output outsig;
  assign outsig = in_0;
endmodule
